// tb.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module tb (
	);

	wire         clock_reset_inst_clock_clk;                                                                   // clock_reset_inst:clock -> [component_dpi_controller_kernel_3mm_inst:clock, irq_mapper:clk, kernel_3mm_inst:clock, main_dpi_controller_inst:clock, stream_source_dpi_bfm_kernel_3mm_A_inst:clock, stream_source_dpi_bfm_kernel_3mm_B_inst:clock, stream_source_dpi_bfm_kernel_3mm_C_inst:clock, stream_source_dpi_bfm_kernel_3mm_D_inst:clock, stream_source_dpi_bfm_kernel_3mm_E_inst:clock, stream_source_dpi_bfm_kernel_3mm_F_inst:clock, stream_source_dpi_bfm_kernel_3mm_G_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                                 // clock_reset_inst:clock2x -> [component_dpi_controller_kernel_3mm_inst:clock2x, main_dpi_controller_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_A_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_B_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_C_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_D_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_E_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_F_inst:clock2x, stream_source_dpi_bfm_kernel_3mm_G_inst:clock2x]
	wire         component_dpi_controller_kernel_3mm_inst_component_call_valid;                                // component_dpi_controller_kernel_3mm_inst:start -> kernel_3mm_inst:start
	wire         kernel_3mm_inst_call_stall;                                                                   // kernel_3mm_inst:busy -> component_dpi_controller_kernel_3mm_inst:busy
	wire         component_dpi_controller_kernel_3mm_inst_component_done_conduit;                              // component_dpi_controller_kernel_3mm_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                                           // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_kernel_3mm_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_kernel_3mm_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_kernel_3mm_inst_dpi_control_bind_conduit;                            // component_dpi_controller_kernel_3mm_inst:bind_interfaces -> kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_kernel_3mm_inst_dpi_control_enable_conduit;                          // component_dpi_controller_kernel_3mm_inst:enable_interfaces -> kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         concatenate_component_done_inst_out_conduit_conduit;                                          // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                        // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         split_component_start_inst_out_conduit_0_conduit;                                             // split_component_start_inst:out_conduit_0 -> component_dpi_controller_kernel_3mm_inst:component_enabled
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_kernel_3mm_A_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_kernel_3mm_A_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_kernel_3mm_A_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_kernel_3mm_B_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_kernel_3mm_B_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_kernel_3mm_B_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_kernel_3mm_C_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_kernel_3mm_C_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_kernel_3mm_C_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_kernel_3mm_D_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_kernel_3mm_D_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_kernel_3mm_D_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_kernel_3mm_E_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_kernel_3mm_E_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_kernel_3mm_E_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_5 -> stream_source_dpi_bfm_kernel_3mm_F_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_5 -> stream_source_dpi_bfm_kernel_3mm_F_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_5 -> stream_source_dpi_bfm_kernel_3mm_F_inst:source_ready
	wire         kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit;           // kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_6 -> stream_source_dpi_bfm_kernel_3mm_G_inst:do_bind
	wire         kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit;         // kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_6 -> stream_source_dpi_bfm_kernel_3mm_G_inst:enable
	wire         kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit; // kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_6 -> stream_source_dpi_bfm_kernel_3mm_G_inst:source_ready
	wire         component_dpi_controller_kernel_3mm_inst_read_implicit_streams_conduit;                       // component_dpi_controller_kernel_3mm_inst:read_implicit_streams -> kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                                  // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         kernel_3mm_inst_return_valid;                                                                 // kernel_3mm_inst:done -> component_dpi_controller_kernel_3mm_inst:done
	wire         component_dpi_controller_kernel_3mm_inst_component_return_stall;                              // component_dpi_controller_kernel_3mm_inst:stall -> kernel_3mm_inst:stall
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_a_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_A_inst:source_data -> kernel_3mm_inst:A
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_b_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_B_inst:source_data -> kernel_3mm_inst:B
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_c_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_C_inst:source_data -> kernel_3mm_inst:C
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_d_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_D_inst:source_data -> kernel_3mm_inst:D
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_e_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_E_inst:source_data -> kernel_3mm_inst:E
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_f_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_F_inst:source_data -> kernel_3mm_inst:F
	wire  [63:0] stream_source_dpi_bfm_kernel_3mm_g_inst_source_data_data;                                     // stream_source_dpi_bfm_kernel_3mm_G_inst:source_data -> kernel_3mm_inst:G
	wire         clock_reset_inst_reset_reset;                                                                 // clock_reset_inst:resetn -> [component_dpi_controller_kernel_3mm_inst:resetn, irq_mapper:reset, kernel_3mm_inst:resetn, main_dpi_controller_inst:resetn, stream_source_dpi_bfm_kernel_3mm_A_inst:resetn, stream_source_dpi_bfm_kernel_3mm_B_inst:resetn, stream_source_dpi_bfm_kernel_3mm_C_inst:resetn, stream_source_dpi_bfm_kernel_3mm_D_inst:resetn, stream_source_dpi_bfm_kernel_3mm_E_inst:resetn, stream_source_dpi_bfm_kernel_3mm_F_inst:resetn, stream_source_dpi_bfm_kernel_3mm_G_inst:resetn]
	wire         component_dpi_controller_kernel_3mm_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_kernel_3mm_inst:done_irq

	clock_reset clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //  output,  width = 1,      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //  output,  width = 1,      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //  output,  width = 1,    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  //   input,  width = 1, reset_ctrl.conduit
	);

	dpic_kernel_3mm component_dpi_controller_kernel_3mm_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                        //   input,   width = 1,                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                      //   input,   width = 1,                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                      //   input,   width = 1,                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_kernel_3mm_inst_dpi_control_bind_conduit),                 //  output,   width = 1,                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_kernel_3mm_inst_dpi_control_enable_conduit),               //  output,   width = 1,               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                  //   input,   width = 1,                component_enabled.conduit
		.component_done                   (component_dpi_controller_kernel_3mm_inst_component_done_conduit),                   //  output,   width = 1,                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_kernel_3mm_inst_component_wait_for_stream_writes_conduit), //  output,   width = 1, component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                                  //   input,   width = 1,                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_kernel_3mm_inst_read_implicit_streams_conduit),            //  output,   width = 1,            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                                  //  output,   width = 1,             readback_from_agents.conduit
		.start                            (component_dpi_controller_kernel_3mm_inst_component_call_valid),                     //  output,   width = 1,                   component_call.valid
		.busy                             (kernel_3mm_inst_call_stall),                                                        //   input,   width = 1,                                 .stall
		.done                             (kernel_3mm_inst_return_valid),                                                      //   input,   width = 1,                 component_return.valid
		.stall                            (component_dpi_controller_kernel_3mm_inst_component_return_stall),                   //  output,   width = 1,                                 .stall
		.done_irq                         (component_dpi_controller_kernel_3mm_inst_component_irq_irq),                        //   input,   width = 1,                    component_irq.irq
		.returndata                       ()                                                                                   //   input,  width = 64,                       returndata.data
	);

	cat_done concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),             //  output,  width = 1,  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_kernel_3mm_inst_component_done_conduit)  //   input,  width = 1, in_conduit_0.conduit
	);

	cat_cwfsw concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),             //  output,  width = 1,  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_kernel_3mm_inst_component_wait_for_stream_writes_conduit)  //   input,  width = 1, in_conduit_0.conduit
	);

	kernel_3mm_cfan kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_kernel_3mm_inst_dpi_control_bind_conduit),                  //   input,  width = 1,    in_conduit.conduit
		.out_conduit_0 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), //  output,  width = 1, out_conduit_0.conduit
		.out_conduit_1 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), //  output,  width = 1, out_conduit_1.conduit
		.out_conduit_2 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), //  output,  width = 1, out_conduit_2.conduit
		.out_conduit_3 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), //  output,  width = 1, out_conduit_3.conduit
		.out_conduit_4 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit), //  output,  width = 1, out_conduit_4.conduit
		.out_conduit_5 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit), //  output,  width = 1, out_conduit_5.conduit
		.out_conduit_6 (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit)  //  output,  width = 1, out_conduit_6.conduit
	);

	kernel_3mm_en_cfan kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_kernel_3mm_inst_dpi_control_enable_conduit),                  //   input,  width = 1,    in_conduit.conduit
		.out_conduit_0 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), //  output,  width = 1, out_conduit_0.conduit
		.out_conduit_1 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), //  output,  width = 1, out_conduit_1.conduit
		.out_conduit_2 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), //  output,  width = 1, out_conduit_2.conduit
		.out_conduit_3 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), //  output,  width = 1, out_conduit_3.conduit
		.out_conduit_4 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit), //  output,  width = 1, out_conduit_4.conduit
		.out_conduit_5 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit), //  output,  width = 1, out_conduit_5.conduit
		.out_conduit_6 (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit)  //  output,  width = 1, out_conduit_6.conduit
	);

	kernel_3mm_ir_cfan kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_kernel_3mm_inst_read_implicit_streams_conduit),                       //   input,  width = 1,    in_conduit.conduit
		.out_conduit_0 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //  output,  width = 1, out_conduit_0.conduit
		.out_conduit_1 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //  output,  width = 1, out_conduit_1.conduit
		.out_conduit_2 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //  output,  width = 1, out_conduit_2.conduit
		.out_conduit_3 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //  output,  width = 1, out_conduit_3.conduit
		.out_conduit_4 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit), //  output,  width = 1, out_conduit_4.conduit
		.out_conduit_5 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit), //  output,  width = 1, out_conduit_5.conduit
		.out_conduit_6 (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit)  //  output,  width = 1, out_conduit_6.conduit
	);

	kernel_3mm kernel_3mm_inst (
		.clock  (clock_reset_inst_clock_clk),                                      //   input,   width = 1,  clock.clk
		.resetn (clock_reset_inst_reset_reset),                                    //   input,   width = 1,  reset.reset_n
		.start  (component_dpi_controller_kernel_3mm_inst_component_call_valid),   //   input,   width = 1,   call.valid
		.busy   (kernel_3mm_inst_call_stall),                                      //  output,   width = 1,       .stall
		.done   (kernel_3mm_inst_return_valid),                                    //  output,   width = 1, return.valid
		.stall  (component_dpi_controller_kernel_3mm_inst_component_return_stall), //   input,   width = 1,       .stall
		.A      (stream_source_dpi_bfm_kernel_3mm_a_inst_source_data_data),        //   input,  width = 64,      A.data
		.B      (stream_source_dpi_bfm_kernel_3mm_b_inst_source_data_data),        //   input,  width = 64,      B.data
		.C      (stream_source_dpi_bfm_kernel_3mm_c_inst_source_data_data),        //   input,  width = 64,      C.data
		.D      (stream_source_dpi_bfm_kernel_3mm_d_inst_source_data_data),        //   input,  width = 64,      D.data
		.E      (stream_source_dpi_bfm_kernel_3mm_e_inst_source_data_data),        //   input,  width = 64,      E.data
		.F      (stream_source_dpi_bfm_kernel_3mm_f_inst_source_data_data),        //   input,  width = 64,      F.data
		.G      (stream_source_dpi_bfm_kernel_3mm_g_inst_source_data_data)         //   input,  width = 64,      G.data
	);

	main_dpi_controller main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //   input,  width = 1,                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //   input,  width = 1,                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //   input,  width = 1,                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //  output,  width = 1,                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //   input,  width = 1,                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), //   input,  width = 1, component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //  output,  width = 1,                       reset_ctrl.conduit
	);

	sp_cstart split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //   input,  width = 1,    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    //  output,  width = 1, out_conduit_0.conduit
	);

	sso_kernel_3mm_A stream_source_dpi_bfm_kernel_3mm_a_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_a_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_B stream_source_dpi_bfm_kernel_3mm_b_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_b_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_C stream_source_dpi_bfm_kernel_3mm_c_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_c_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_D stream_source_dpi_bfm_kernel_3mm_d_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_d_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_3_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_E stream_source_dpi_bfm_kernel_3mm_e_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_e_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_4_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_F stream_source_dpi_bfm_kernel_3mm_f_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_5_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_5_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_f_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_5_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	sso_kernel_3mm_G stream_source_dpi_bfm_kernel_3mm_g_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                   //   input,   width = 1,              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                 //   input,   width = 1,              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                 //   input,   width = 1,            clock2x.clk
		.do_bind      (kernel_3mm_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_6_conduit),           //   input,   width = 1,   dpi_control_bind.conduit
		.enable       (kernel_3mm_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_6_conduit),         //   input,   width = 1, dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_kernel_3mm_g_inst_source_data_data),                                     //  output,  width = 64,        source_data.data
		.source_ready (kernel_3mm_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_6_conduit), //   input,   width = 1,       source_ready.conduit
		.source_valid ()                                                                                              //  output,   width = 1,             source.conduit
	);

	tb_altera_irq_mapper_1920_trjgw7i irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                                 //   input,  width = 1,       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                              //   input,  width = 1, clk_reset.reset
		.sender_irq (component_dpi_controller_kernel_3mm_inst_component_irq_irq)  //  output,  width = 1,    sender.irq
	);

endmodule
