    .INIT_00(256'h022ffd207311d800022ffd2073119801022ffd2500036218022ffd206e31e010),
    .INIT_01(256'h022ffd2073101004022ffd2073120ab4022ffd20731221e5022ffd2073132206),
    .INIT_02(256'h022ffd0b0320b032022ffd250002f013022ffd207310b002022ffd207312f01f),
    .INIT_03(256'h022ffd2071f20793022ffd20707206e3022ffd368123220f022ffd1d0001d002),
    .INIT_04(256'h022ffd207071d002022ffd25000324f8022ffd206e31d001022ffd207250b032),
    .INIT_05(256'h022ffd2500022008022ffd206e320754022ffd2070301004022ffd20719324f8),
    .INIT_06(256'h022ffd2070b0b016022ffd3681f2f03a022ffd1d00011001022ffd0b0320b03a),
    .INIT_07(256'h022ffd250000b018022ffd206e31f000022ffd207090b017022ffd2071d1d000),
    .INIT_08(256'h022ffd206e30b01a022ffd207071f000022ffd207070b019022ffd2070b1f000),
    .INIT_09(256'h022ffd206e50b01c022ffd207031f000022ffd207210b01b022ffd207f01f000),
    .INIT_0A(256'h022ffd0401036017022ffd0b00f1f000022ffd141060b01d022ffd0b1131f000),
    .INIT_0B(256'h022ffd206ce32481022ffd206c41d001022ffd206c40b032022ffd00c00208ac),
    .INIT_0C(256'h022ffd0b00d01001022ffd206bc22008022ffd0b00e324d4022ffd207371d002),
    .INIT_0D(256'h022ffd206e30bf12022ffd206bc0be11022ffd0b00c0bd10022ffd206bc2f01e),
    .INIT_0E(256'h022ffd206ef2fd10022ffd206e513f00022ffd2070313e00022ffd2071911d01),
    .INIT_0F(256'h022ffd0401020b66022ffd0b0122ff12022ffd1410603f01022ffd0b1132fe11),
    .INIT_10(256'h022ffd0b0100b03b022ffd206bc2f00f022ffd0b01103001022ffd206bc0b00f),
    .INIT_11(256'h022ffd0bc171c0e0022ffd2500003e7e022ffd206e30be0e022ffd206bc0307e),
    .INIT_12(256'h022ffd1dcff0b016022ffd0bc1620918022ffd3488520901022ffd1dcff36264),
    .INIT_13(256'h022ffd348850b018022ffd1dcff1f000022ffd0bc190b017022ffd3488b1d000),
    .INIT_14(256'h022ffd0bc1b0b01a022ffd3488b1f000022ffd1dcff0b019022ffd0bc181f000),
    .INIT_15(256'h022ffd1dcff0b01c022ffd0bc1a1f000022ffd348850b01b022ffd1dcff1f000),
    .INIT_16(256'h022ffd348853625d022ffd1dcff1f000022ffd0bc1d0b01d022ffd3488b1f000),
    .INIT_17(256'h022ffd25000206e3022ffd3488b20782022ffd1dcff20763022ffd0bc1c22264),
    .INIT_18(256'h022ffd0bc1722008022ffd3286920754022ffd1dd0001004022ffd0bd2020793),
    .INIT_19(256'h022ffd0bc202b80f022ffd208912b40f022ffd0bc162b20f022ffd20885208ac),
    .INIT_1A(256'h022ffd3287222008022ffd1dd0020782022ffd0bd2120754022ffd2089701002),
    .INIT_1B(256'h022ffd208910d004022ffd0bc180900e022ffd208852f032022ffd0bc1901000),
    .INIT_1C(256'h022ffd1dd0009018022ffd0bd222f007022ffd2089709017022ffd0bc213229d),
    .INIT_1D(256'h022ffd0bc1a0901a022ffd208852f009022ffd0bc1b09019022ffd3287b2f008),
    .INIT_1E(256'h022ffd0bd232b04e022ffd208972f00b022ffd0bc220901b022ffd208912f00a),
    .INIT_1F(256'h022ffd2088509002022ffd0bc1d36283022ffd328841d0a0022ffd1dd00030f0),
    .INIT_20(256'h022ffd208971d0e0022ffd0bc23223f6022ffd20891323f5022ffd0bc1c0d002),
    .INIT_21(256'h022ffd206e536290022ffd207091d0b0022ffd2072f223f5022ffd2500036286),
    .INIT_22(256'h022ffd2070520725022ffd250002dc01022ffd206e503c0f022ffd206bd0bc07),
    .INIT_23(256'h022ffd206e322003022ffd206bd206e3022ffd206e5206bd022ffd20729206e5),
    .INIT_24(256'h022ffd206e522412022ffd207292072b022ffd2070536294022ffd250001d0d0),
    .INIT_25(256'h022ffd2071922402022ffd2500020709022ffd206e536298022ffd206bd1d0f0),
    .INIT_26(256'h022ffd206e33241b022ffd206bd0d080022ffd206e53241b022ffd2072d1d0c0),
    .INIT_27(256'h022ffd2b1bb363f5022ffd2b00a0d020022ffd2b0090900d022ffd25000223f3),
    .INIT_28(256'h022ffd208b509002022ffd01c00362a7022ffd209101d04f022ffd2b08e09006),
    .INIT_29(256'h022ffd208b51d053022ffd01c10223f6022ffd25000323f5022ffd200590d002),
    .INIT_2A(256'h022ffd250002078b022ffd208b5206e3022ffd01c0720727022ffd25000362ae),
    .INIT_2B(256'h022ffd01c01362c5022ffd250001d052022ffd208b5223f4022ffd01c0d2079a),
    .INIT_2C(256'h022ffd208b51d020022ffd01c0409006022ffd250002073a022ffd208b520725),
    .INIT_2D(256'h022ffd01f0009006022ffd01e002073a022ffd01d00206e5022ffd25000363f3),
    .INIT_2E(256'h022ffd208db2073a022ffd01100206ef022ffd01080363f3022ffd208e41d030),
    .INIT_2F(256'h022ffd2b00a2d001022ffd2b3893a3f3022ffd25000206b0022ffd208c409006),
    .INIT_30(256'h022ffd25000206e3022ffd2091020737022ffd2b08e206ce022ffd2b63b00100),
    .INIT_31(256'h022ffd2b08e2072b022ffd2b37b362c9022ffd2b00a1d055022ffd2b1c922003),
    .INIT_32(256'h022ffd2b72a20709022ffd2b649362cd022ffd250001d044022ffd2091022412),
    .INIT_33(256'h022ffd250002071d022ffd20910362de022ffd2b08e1d04e022ffd2b0bb22402),
    .INIT_34(256'h022ffd2b08e363f3022ffd2b57b1d020022ffd2b20a09006022ffd2b6492073a),
    .INIT_35(256'h022ffd2b63b3a3f3022ffd2b20a206d3022ffd2b6c90120a022ffd20910206e5),
    .INIT_36(256'h022ffd2b00a2fd0a022ffd250002fc09022ffd209102fb08022ffd2b08e2fa07),
    .INIT_37(256'h022ffd2b00a36331022ffd2d1081d054022ffd2d00822427022ffd2b4192fe0b),
    .INIT_38(256'h022ffd250001d020022ffd2d10809006022ffd2d0082073a022ffd2b25920729),
    .INIT_39(256'h022ffd2dd08206d3022ffd2dc080120a022ffd2b289206e5022ffd2b00a363f3),
    .INIT_3A(256'h022ffd2b00a1dec0022ffd250002fb3f022ffd2df082fa3e022ffd2de083a3f3),
    .INIT_3B(256'h022ffd09e08223f3022ffd09d08322f0022ffd09c080de80022ffd2b2893230f),
    .INIT_3C(256'h022ffd208eb0ba02022ffd208be206a9022ffd25000206a9022ffd09f08206a9),
    .INIT_3D(256'h022ffd250002fc0c022ffd208c4206a9022ffd208e4363f3022ffd2500018fa0),
    .INIT_3E(256'h022ffd0bf0f20ab4022ffd208db2ff0f022ffd011002fe0e022ffd010202fd0d),
    .INIT_3F(256'h022ffd208f50bf12022ffd0bc0c0be11022ffd0bd0d0bd10022ffd0be0e206e3),
    .INIT_40(256'h022ffd208ca00ce0022ffd208b2206bd022ffd208f800cf0022ffd2500020707),
    .INIT_41(256'h022ffd208f80bc3f022ffd25000206bd022ffd2090700cd0022ffd25000206bd),
    .INIT_42(256'h022ffd208be20737022ffd208db206ce022ffd01101206c4022ffd01080206c4),
    .INIT_43(256'h022ffd25000206a9022ffd208d0223f3022ffd208af206bd022ffd208c40bc3e),
    .INIT_44(256'h022ffd2500018ea0022ffd369100ba02022ffd0d008206a9022ffd0900e206a9),
    .INIT_45(256'h022ffd250002fd11022ffd329142fc10022ffd0d002206a9022ffd0900e363f3),
    .INIT_46(256'h022ffd2f1170bf0c022ffd2f116206e3022ffd0110020b66022ffd370012fe12),
    .INIT_47(256'h022ffd2f11b206c4022ffd2f11a0bc0f022ffd2f1190bd0e022ffd2f1180be0d),
    .INIT_48(256'h022ffd2b6c900cd0022ffd0108420737022ffd2f11d206ce022ffd2f11c206c4),
    .INIT_49(256'h022ffd2092e00cf0022ffd11001206bd022ffd2b00b00ce0022ffd2b00a206bd),
    .INIT_4A(256'h022ffd36926206c4022ffd1d0ff206c4022ffd2098d0bc3f022ffd20933206bd),
    .INIT_4B(256'h022ffd09d08206bd022ffd09c080bc3e022ffd2500020737022ffd37000206ce),
    .INIT_4C(256'h022ffd1d0c109002022ffd250003634f022ffd09f081d058022ffd09e08223f3),
    .INIT_4D(256'h022ffd001f02073a022ffd3295e20731022ffd1d0c23e34f022ffd329490d004),
    .INIT_4E(256'h022ffd001d0206e5022ffd2097c363f3022ffd001e01d020022ffd2097c09006),
    .INIT_4F(256'h022ffd01100206e3022ffd2097c3a3f3022ffd001c0206d3022ffd2097c01208),
    .INIT_50(256'h022ffd2f12e2fd3b022ffd2f12c2fc36022ffd2f12a2fb35022ffd2f1282fa34),
    .INIT_51(256'h022ffd2f12f0bf3b022ffd2f12d0be36022ffd2f12b0bd35022ffd2f1290bc34),
    .INIT_52(256'h022ffd001e02062f022ffd2097c20681022ffd001f001b00022ffd2500001a01),
    .INIT_53(256'h022ffd001c01d051022ffd2097c223f3022ffd001d0206bd022ffd2097c09c07),
    .INIT_54(256'h022ffd2f52c09006022ffd2f62a2073a022ffd2f72820723022ffd2097c36397),
    .INIT_55(256'h022ffd016000120a022ffd01500206e5022ffd01400363f3022ffd2f42e1d020),
    .INIT_56(256'h022ffd2f52d3236b022ffd2f62b1dec0022ffd2f7293a3f3022ffd01700206d3),
    .INIT_57(256'h022ffd2097c206a9022ffd001f0223f3022ffd229483235f022ffd2f42f0de80),
    .INIT_58(256'h022ffd2097c18fa0022ffd001d00ba02022ffd2097c206a9022ffd001e0206a9),
    .INIT_59(256'h022ffd0310f2fd0d022ffd001702fc0c022ffd2097c206a9022ffd001c0363f3),
    .INIT_5A(256'h022ffd0310f206a9022ffd0016022381022ffd037f02ff0f022ffd2f1292fe0e),
    .INIT_5B(256'h022ffd0310f18ea0022ffd001500ba02022ffd036f0206a9022ffd2f12b206a9),
    .INIT_5C(256'h022ffd0310f2fd11022ffd001402fc10022ffd035f0206a9022ffd2f12d363f3),
    .INIT_5D(256'h022ffd2f1280b206022ffd011000b105022ffd034f00b004022ffd2f12f2fe12),
    .INIT_5E(256'h022ffd229483e3f3022ffd2f12e1ae20022ffd2f12c1ad10022ffd2f12a18c00),
    .INIT_5F(256'h022ffd145002f40f022ffd1410003401022ffd144000b40f022ffd1410020b66),
    .INIT_60(256'h022ffd14700206e3022ffd1410020901022ffd146002089d022ffd1410022381),
    .INIT_61(256'h022ffd1450009f08022ffd141000127b022ffd144002b6c9022ffd141002b00a),
    .INIT_62(256'h022ffd14700206bd022ffd1410009c08022ffd1460009d08022ffd1410009e08),
    .INIT_63(256'h022ffd0b929206bd022ffd0b82800ce0022ffd00170206bd022ffd2500000cd0),
    .INIT_64(256'h022ffd01b0019201022ffd20a58206e3022ffd20a3a206bd022ffd20a2e00cf0),
    .INIT_65(256'h022ffd0ba261d050022ffd14b00223f4022ffd14a0e208ac022ffd0ba2536387),
    .INIT_66(256'h022ffd14b0009006022ffd14a002073a022ffd14b0020721022ffd14a00363f5),
    .INIT_67(256'h022ffd062b001202022ffd0b217206e5022ffd14b00363f3022ffd14a001d020),
    .INIT_68(256'h022ffd14a00206a9022ffd14b00206a9022ffd14a003a3f3022ffd2f217206d3),
    .INIT_69(256'h022ffd14a00363f3022ffd14b0018bc0022ffd14a000bc02022ffd14b00206a9),
    .INIT_6A(256'h022ffd0ba270d040022ffd14b0009002022ffd14a00206a9022ffd14b00206a9),
    .INIT_6B(256'h022ffd14b00323e1022ffd14a001fb00022ffd14b001da00022ffd14a00363e1),
    .INIT_6C(256'h022ffd06b201da80022ffd0b216323e1022ffd14b001fb00022ffd14a001da20),
    .INIT_6D(256'h022ffd0b92b1fb00022ffd0b82a1daa0022ffd00160323e1022ffd2fb161fb00),
    .INIT_6E(256'h022ffd01b00323e1022ffd20a581fb00022ffd20a3a1dac0022ffd20a2e323e1),
    .INIT_6F(256'h022ffd0ba261da20022ffd14b00323e1022ffd14a0e1fb00022ffd0ba251dae0),
    .INIT_70(256'h022ffd14b001fb01022ffd14a001da80022ffd14b00323e1022ffd14a001fb01),
    .INIT_71(256'h022ffd062b0323e1022ffd0b2191fb01022ffd14b001daa0022ffd14a00323e1),
    .INIT_72(256'h022ffd14a001da00022ffd14b00323e1022ffd14a001fb01022ffd2f2191dac0),
    .INIT_73(256'h022ffd14a001fb02022ffd14b001da20022ffd14a00323e1022ffd14b001fb02),
    .INIT_74(256'h022ffd0ba27323e1022ffd14b001fb02022ffd14a001da80022ffd14b00323e1),
    .INIT_75(256'h022ffd14b001dac0022ffd14a00323e1022ffd14b001fb02022ffd14a001daa0),
    .INIT_76(256'h022ffd06b201fb03022ffd0b2181da00022ffd14b00323e1022ffd14a001fb02),
    .INIT_77(256'h022ffd0b92d323e1022ffd0b82c1fb03022ffd001501dae0022ffd2fb18323e1),
    .INIT_78(256'h022ffd01b00000a0022ffd20a582089d022ffd20a3a206e3022ffd20a2e223f3),
    .INIT_79(256'h022ffd0ba26208eb022ffd14b00208be022ffd14a0e208db022ffd0ba25001b0),
    .INIT_7A(256'h022ffd14b0000ce0022ffd14a00206bd022ffd14b0000cf0022ffd14a0000bc0),
    .INIT_7B(256'h022ffd062b000cb0022ffd0b21b206bd022ffd14b0000cd0022ffd14a00206bd),
    .INIT_7C(256'h022ffd14a00206e3022ffd14b00223f3022ffd14a00208ac022ffd2f21b206bd),
    .INIT_7D(256'h022ffd14a00206e3022ffd14b002071f022ffd14a0022008022ffd14b0020782),
    .INIT_7E(256'h022ffd0ba272b20f022ffd14b00208ac022ffd14a002013e022ffd14b002089d),
    .INIT_7F(256'h022ffd14b002075402bff314a000100202bff014b002b80f022ffd14a002b40f),
    .INITP_00(256'h61ff4d575571d1f3f8f6c2d04ae56f5cd1d7e756f463dd55d8cd4d53584ffde4),
    .INITP_01(256'he97fe04d65e4515a6c5873cc765573cb7fed795b61eae0d6f2c04ec376dc535d),
    .INITP_02(256'h66fdcb6d7d41e5f9cb71e941e2f9ceeaef417bea49637d5866e6695bf4c67ac5),
    .INITP_03(256'h75786df34ee474e0eb64f77cff4ffc61607f6674e8e4c665f5fe6cf67ff6e2db),
    .INITP_04(256'h484fd27e7c53fb51c0e4644d695fda706bd1f5d1c56276c6635a4efc7a61e576),
    .INITP_05(256'hd174e248c8c15bd57e4340fc79e5e162ed79737aedebf17177e36bdbf4f3e7ec),
    .INITP_06(256'h53eecd6ad0766ce0ca6ccb70ef65f6edeb6c6261f4faf369f86054f566f6fdc1),
    .INITP_07(256'hd2f0495c795fdee7735854635d7eefd96bf1454744fa476df2d14f51f46b56d9),
    .INITP_08(256'h4f4f405fd1dedae9f57172c96eca74daef4bf54172c750cbc2e07de0c5f056e0),
    .INITP_09(256'h4057e7ca79d669d5e24dd240cdf2cd6b7247e3ed5543c76b6f54df4dc5584ad2),
    .INITP_0A(256'hc57df04c6ae9c5c2e166dc56e5fb4ed1fd54fc48fd4878f54eda584d59cdc0d5),
    .INITP_0B(256'hc2f5e2fff655cedec1c1634e7b5bc6d9e04b414d61ccfbc173d2c57e49e9c572),
    .INITP_0C(256'hc6457d567e43e85d617f426ec3c86be8fa4b416b62e649e8c0edfff9e4f0dbf0),
    .INITP_0D(256'hf6e547f0c051ed6d7e5f5bc5f05e7ec9e55d6052e4f84d6e5eecd66e4d6edf40),
    .INITP_0E(256'h62c6524464c1e5d8e7c6fb45e3fbcfe5d8eac6fb43e5de59c04666c6fdcfe5de),
    .INITP_0F(256'he578c6d2767b44fbc4ef5ae8c4ff58444e41ea42e94260ccec77cae5d9d4ed77),
