library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;
use std.textio.all;

use work.sim_package.all;



entity bicg_tb is

end entity bicg_tb;

architecture behav of bicg_tb is

	-- Constant declarations

	constant HALF_CLK_PERIOD : TIME := 2.00 ns;
	constant TRANSACTION_NUM : INTEGER := 1;
	constant INPUT_end : STRING := "";
	constant OUTPUT_end : STRING := "../VHDL_OUT/output_end.dat";
	constant DATA_WIDTH_end : INTEGER := 32;
	constant INPUT_A : STRING := "../INPUT_VECTORS/input_A.dat";
	constant OUTPUT_A : STRING := "";
	constant DATA_WIDTH_A : INTEGER := 32;
	constant ADDR_WIDTH_A : INTEGER := 32;
	constant DATA_DEPTH_A : INTEGER := 900;
	constant INPUT_s : STRING := "../INPUT_VECTORS/input_s.dat";
	constant OUTPUT_s : STRING := "../VHDL_OUT/output_s.dat";
	constant DATA_WIDTH_s : INTEGER := 32;
	constant ADDR_WIDTH_s : INTEGER := 32;
	constant DATA_DEPTH_s : INTEGER := 30;
	constant INPUT_q : STRING := "../INPUT_VECTORS/input_q.dat";
	constant OUTPUT_q : STRING := "../VHDL_OUT/output_q.dat";
	constant DATA_WIDTH_q : INTEGER := 32;
	constant ADDR_WIDTH_q : INTEGER := 32;
	constant DATA_DEPTH_q : INTEGER := 30;
	constant INPUT_p : STRING := "../INPUT_VECTORS/input_p.dat";
	constant OUTPUT_p : STRING := "";
	constant DATA_WIDTH_p : INTEGER := 32;
	constant ADDR_WIDTH_p : INTEGER := 32;
	constant DATA_DEPTH_p : INTEGER := 30;
	constant INPUT_r : STRING := "../INPUT_VECTORS/input_r.dat";
	constant OUTPUT_r : STRING := "";
	constant DATA_WIDTH_r : INTEGER := 32;
	constant ADDR_WIDTH_r : INTEGER := 32;
	constant DATA_DEPTH_r : INTEGER := 30;

	-- Signal declarations

	signal tb_clk : std_logic := '0';
	signal tb_rst : std_logic := '0';
	signal tb_start_valid : std_logic := '0';
	signal tb_start_ready : std_logic;
	signal tb_end_valid : std_logic;

	signal end_mem_ce0 : std_logic;
	signal end_mem_we0 : std_logic;
	signal end_mem_dout0 : std_logic_vector(DATA_WIDTH_end - 1 downto 0);
	signal end_mem_din0 : std_logic_vector(DATA_WIDTH_end - 1 downto 0);


	signal A_mem_ce0 : std_logic;
	signal A_mem_we0 : std_logic;
	signal A_mem_din0 : std_logic_vector(DATA_WIDTH_A - 1 downto 0);
	signal A_mem_dout0 : std_logic_vector(DATA_WIDTH_A - 1 downto 0);
	signal A_mem_address0 : std_logic_vector(ADDR_WIDTH_A - 1 downto 0);

	signal A_mem_ce1 : std_logic;
	signal A_mem_we1 : std_logic;
	signal A_mem_din1 : std_logic_vector(DATA_WIDTH_A - 1 downto 0);
	signal A_mem_dout1 : std_logic_vector(DATA_WIDTH_A - 1 downto 0);
	signal A_mem_address1 : std_logic_vector(ADDR_WIDTH_A - 1 downto 0);

	signal s_mem_ce0 : std_logic;
	signal s_mem_we0 : std_logic;
	signal s_mem_din0 : std_logic_vector(DATA_WIDTH_s - 1 downto 0);
	signal s_mem_dout0 : std_logic_vector(DATA_WIDTH_s - 1 downto 0);
	signal s_mem_address0 : std_logic_vector(ADDR_WIDTH_s - 1 downto 0);

	signal s_mem_ce1 : std_logic;
	signal s_mem_we1 : std_logic;
	signal s_mem_din1 : std_logic_vector(DATA_WIDTH_s - 1 downto 0);
	signal s_mem_dout1 : std_logic_vector(DATA_WIDTH_s - 1 downto 0);
	signal s_mem_address1 : std_logic_vector(ADDR_WIDTH_s - 1 downto 0);

	signal q_mem_ce0 : std_logic;
	signal q_mem_we0 : std_logic;
	signal q_mem_din0 : std_logic_vector(DATA_WIDTH_q - 1 downto 0);
	signal q_mem_dout0 : std_logic_vector(DATA_WIDTH_q - 1 downto 0);
	signal q_mem_address0 : std_logic_vector(ADDR_WIDTH_q - 1 downto 0);

	signal q_mem_ce1 : std_logic;
	signal q_mem_we1 : std_logic;
	signal q_mem_din1 : std_logic_vector(DATA_WIDTH_q - 1 downto 0);
	signal q_mem_dout1 : std_logic_vector(DATA_WIDTH_q - 1 downto 0);
	signal q_mem_address1 : std_logic_vector(ADDR_WIDTH_q - 1 downto 0);

	signal p_mem_ce0 : std_logic;
	signal p_mem_we0 : std_logic;
	signal p_mem_din0 : std_logic_vector(DATA_WIDTH_p - 1 downto 0);
	signal p_mem_dout0 : std_logic_vector(DATA_WIDTH_p - 1 downto 0);
	signal p_mem_address0 : std_logic_vector(ADDR_WIDTH_p - 1 downto 0);

	signal p_mem_ce1 : std_logic;
	signal p_mem_we1 : std_logic;
	signal p_mem_din1 : std_logic_vector(DATA_WIDTH_p - 1 downto 0);
	signal p_mem_dout1 : std_logic_vector(DATA_WIDTH_p - 1 downto 0);
	signal p_mem_address1 : std_logic_vector(ADDR_WIDTH_p - 1 downto 0);

	signal r_mem_ce0 : std_logic;
	signal r_mem_we0 : std_logic;
	signal r_mem_din0 : std_logic_vector(DATA_WIDTH_r - 1 downto 0);
	signal r_mem_dout0 : std_logic_vector(DATA_WIDTH_r - 1 downto 0);
	signal r_mem_address0 : std_logic_vector(ADDR_WIDTH_r - 1 downto 0);

	signal r_mem_ce1 : std_logic;
	signal r_mem_we1 : std_logic;
	signal r_mem_din1 : std_logic_vector(DATA_WIDTH_r - 1 downto 0);
	signal r_mem_dout1 : std_logic_vector(DATA_WIDTH_r - 1 downto 0);
	signal r_mem_address1 : std_logic_vector(ADDR_WIDTH_r - 1 downto 0);


	signal tb_temp_idle : std_logic:= '1';
	shared variable transaction_idx : INTEGER := 0;

begin


duv: 	 entity work.bicg
		port map (
			clk => tb_clk,
			rst => tb_rst,
			end_out => end_mem_din0,
			end_valid => tb_end_valid,
			end_ready => '1',
			A_address0 => A_mem_address0,
			A_ce0 => A_mem_ce0,
			A_we0 => A_mem_we0,
			A_din0 => A_mem_dout0,
			A_dout0 => A_mem_din0,
			A_address1 => A_mem_address1,
			A_ce1 => A_mem_ce1,
			A_we1 => A_mem_we1,
			A_din1 => A_mem_dout1,
			A_dout1 => A_mem_din1,
			s_address0 => s_mem_address0,
			s_ce0 => s_mem_ce0,
			s_we0 => s_mem_we0,
			s_din0 => s_mem_dout0,
			s_dout0 => s_mem_din0,
			s_address1 => s_mem_address1,
			s_ce1 => s_mem_ce1,
			s_we1 => s_mem_we1,
			s_din1 => s_mem_dout1,
			s_dout1 => s_mem_din1,
			q_address0 => q_mem_address0,
			q_ce0 => q_mem_ce0,
			q_we0 => q_mem_we0,
			q_din0 => q_mem_dout0,
			q_dout0 => q_mem_din0,
			q_address1 => q_mem_address1,
			q_ce1 => q_mem_ce1,
			q_we1 => q_mem_we1,
			q_din1 => q_mem_dout1,
			q_dout1 => q_mem_din1,
			p_address0 => p_mem_address0,
			p_ce0 => p_mem_ce0,
			p_we0 => p_mem_we0,
			p_din0 => p_mem_dout0,
			p_dout0 => p_mem_din0,
			p_address1 => p_mem_address1,
			p_ce1 => p_mem_ce1,
			p_we1 => p_mem_we1,
			p_din1 => p_mem_dout1,
			p_dout1 => p_mem_din1,
			r_address0 => r_mem_address0,
			r_ce0 => r_mem_ce0,
			r_we0 => r_mem_we0,
			r_din0 => r_mem_dout0,
			r_dout0 => r_mem_din0,
			r_address1 => r_mem_address1,
			r_ce1 => r_mem_ce1,
			r_we1 => r_mem_we1,
			r_din1 => r_mem_dout1,
			r_dout1 => r_mem_din1,
			start_in => (others => '0'),
			start_ready => tb_start_ready,
			start_valid => tb_start_valid
		);


arg_inst_end:	 entity work.single_argument
	generic map(
		TV_IN => INPUT_end,
		TV_OUT => OUTPUT_end,
		DATA_WIDTH => DATA_WIDTH_end
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => '1',
		we0 => tb_end_valid,
		mem_dout0 => end_mem_dout0,
		mem_din0 => end_mem_din0,
		done => tb_temp_idle
	);

mem_inst_A:	 entity work.two_port_RAM 
	generic map(
		TV_IN => INPUT_A,
		TV_OUT => OUTPUT_A,
		DEPTH => DATA_DEPTH_A,
		DATA_WIDTH => DATA_WIDTH_A,
		ADDR_WIDTH => ADDR_WIDTH_A
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => A_mem_ce0,
		we0 => A_mem_we0,
		address0 => A_mem_address0,
		mem_dout0 => A_mem_dout0,
		mem_din0 => A_mem_din0,
		ce1 => A_mem_ce1,
		we1 => A_mem_we1,
		address1 => A_mem_address1,
		mem_dout1 => A_mem_dout1,
		mem_din1 => A_mem_din1,
		done => tb_temp_idle
	);

mem_inst_s:	 entity work.two_port_RAM 
	generic map(
		TV_IN => INPUT_s,
		TV_OUT => OUTPUT_s,
		DEPTH => DATA_DEPTH_s,
		DATA_WIDTH => DATA_WIDTH_s,
		ADDR_WIDTH => ADDR_WIDTH_s
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => s_mem_ce0,
		we0 => s_mem_we0,
		address0 => s_mem_address0,
		mem_dout0 => s_mem_dout0,
		mem_din0 => s_mem_din0,
		ce1 => s_mem_ce1,
		we1 => s_mem_we1,
		address1 => s_mem_address1,
		mem_dout1 => s_mem_dout1,
		mem_din1 => s_mem_din1,
		done => tb_temp_idle
	);

mem_inst_q:	 entity work.two_port_RAM 
	generic map(
		TV_IN => INPUT_q,
		TV_OUT => OUTPUT_q,
		DEPTH => DATA_DEPTH_q,
		DATA_WIDTH => DATA_WIDTH_q,
		ADDR_WIDTH => ADDR_WIDTH_q
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => q_mem_ce0,
		we0 => q_mem_we0,
		address0 => q_mem_address0,
		mem_dout0 => q_mem_dout0,
		mem_din0 => q_mem_din0,
		ce1 => q_mem_ce1,
		we1 => q_mem_we1,
		address1 => q_mem_address1,
		mem_dout1 => q_mem_dout1,
		mem_din1 => q_mem_din1,
		done => tb_temp_idle
	);

mem_inst_p:	 entity work.two_port_RAM 
	generic map(
		TV_IN => INPUT_p,
		TV_OUT => OUTPUT_p,
		DEPTH => DATA_DEPTH_p,
		DATA_WIDTH => DATA_WIDTH_p,
		ADDR_WIDTH => ADDR_WIDTH_p
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => p_mem_ce0,
		we0 => p_mem_we0,
		address0 => p_mem_address0,
		mem_dout0 => p_mem_dout0,
		mem_din0 => p_mem_din0,
		ce1 => p_mem_ce1,
		we1 => p_mem_we1,
		address1 => p_mem_address1,
		mem_dout1 => p_mem_dout1,
		mem_din1 => p_mem_din1,
		done => tb_temp_idle
	);

mem_inst_r:	 entity work.two_port_RAM 
	generic map(
		TV_IN => INPUT_r,
		TV_OUT => OUTPUT_r,
		DEPTH => DATA_DEPTH_r,
		DATA_WIDTH => DATA_WIDTH_r,
		ADDR_WIDTH => ADDR_WIDTH_r
	)
	port map(
		clk => tb_clk,
		rst => tb_rst,
		ce0 => r_mem_ce0,
		we0 => r_mem_we0,
		address0 => r_mem_address0,
		mem_dout0 => r_mem_dout0,
		mem_din0 => r_mem_din0,
		ce1 => r_mem_ce1,
		we1 => r_mem_we1,
		address1 => r_mem_address1,
		mem_dout1 => r_mem_dout1,
		mem_din1 => r_mem_din1,
		done => tb_temp_idle
	);



----------------------------------------------------------------------------
-- Write "[[[runtime]]]" and "[[[/runtime]]]" for output transactor
write_output_transactor_end_runtime_proc : process
	file fp             : TEXT;
	variable fstatus    : FILE_OPEN_STATUS;
	variable token_line : LINE;
	variable token      : STRING(1 to 1024);

begin
	file_open(fstatus, fp, OUTPUT_end, WRITE_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_end & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	while transaction_idx /= TRANSACTION_NUM loop
		wait until tb_clk'event and tb_clk = '1';
	end loop;
	wait until tb_clk'event and tb_clk = '1';
	wait until tb_clk'event and tb_clk = '1';
	file_open(fstatus, fp, OUTPUT_end, APPEND_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_end & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[/runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	wait;
end process;
write_output_transactor_s_runtime_proc : process
	file fp             : TEXT;
	variable fstatus    : FILE_OPEN_STATUS;
	variable token_line : LINE;
	variable token      : STRING(1 to 1024);

begin
	file_open(fstatus, fp, OUTPUT_s, WRITE_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_s & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	while transaction_idx /= TRANSACTION_NUM loop
		wait until tb_clk'event and tb_clk = '1';
	end loop;
	wait until tb_clk'event and tb_clk = '1';
	wait until tb_clk'event and tb_clk = '1';
	file_open(fstatus, fp, OUTPUT_s, APPEND_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_s & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[/runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	wait;
end process;
write_output_transactor_q_runtime_proc : process
	file fp             : TEXT;
	variable fstatus    : FILE_OPEN_STATUS;
	variable token_line : LINE;
	variable token      : STRING(1 to 1024);

begin
	file_open(fstatus, fp, OUTPUT_q, WRITE_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_q & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	while transaction_idx /= TRANSACTION_NUM loop
		wait until tb_clk'event and tb_clk = '1';
	end loop;
	wait until tb_clk'event and tb_clk = '1';
	wait until tb_clk'event and tb_clk = '1';
	file_open(fstatus, fp, OUTPUT_q, APPEND_MODE);
	if (fstatus /= OPEN_OK) then
		assert false report "Open file " & OUTPUT_q & " failed!!!" severity note;
		assert false report "ERROR: Simulation using HLS TB failed." severity failure;
	end if;
	write(token_line, string'("[[[/runtime]]]"));
	writeline(fp, token_line);
	file_close(fp);
	wait;
end process;
----------------------------------------------------------------------------



----------------------------------------------------------------------------
generate_sim_done_proc : process
begin
	while (transaction_idx /= TRANSACTION_NUM) loop
		wait until tb_clk'event and tb_clk = '1';
	end loop;
	wait until tb_clk'event and tb_clk = '1';
	wait until tb_clk'event and tb_clk = '1';
	wait until tb_clk'event and tb_clk = '1';
	assert false report "simulation done!" severity note;
	assert false report "NORMAL EXIT (note: failure is to force the simulator to stop)" severity failure;
	wait;
end process;

----------------------------------------------------------------------------
gen_clock_proc : process
begin
	tb_clk <= '0';
	while (true) loop
		wait for HALF_CLK_PERIOD;
		tb_clk <= not tb_clk;
	end loop;
	wait;
end process;

----------------------------------------------------------------------------
gen_reset_proc : process
begin
	tb_rst <= '1';
	wait for 10 ns;
	tb_rst <= '0';
	wait;
end process;

----------------------------------------------------------------------------
generate_idle_signal: process(tb_clk,tb_rst)
begin
   if (tb_rst = '1') then
       tb_temp_idle <= '1';
   elsif rising_edge(tb_clk) then
       tb_temp_idle <= tb_temp_idle;
       if (tb_start_valid = '1') then
           tb_temp_idle <= '0';
       elsif(tb_end_valid = '1') then
           tb_temp_idle <= '1';
       end if;
   end if;
end process generate_idle_signal;

----------------------------------------------------------------------------
generate_start_signal : process(tb_clk, tb_rst)
begin
   if (tb_rst = '1') then
       tb_start_valid <= '0';
   elsif rising_edge(tb_clk) then
       if (tb_temp_idle = '1' and tb_start_ready = '1' and tb_start_valid = '0') then
           tb_start_valid <= '1';
       else
           tb_start_valid <= '0';
       end if;
   end if;
end process generate_start_signal;

----------------------------------------------------------------------------
transaction_increment : process
begin
	wait until tb_rst = '0';
	while (tb_temp_idle /= '1') loop
		wait until tb_clk'event and tb_clk = '1';
	end loop;
	wait until tb_temp_idle = '0';

	while (true) loop
		while (tb_temp_idle /= '1') loop
			wait until tb_clk'event and tb_clk = '1';
		end loop;
		transaction_idx := transaction_idx + 1;
		wait until tb_temp_idle = '0';
	end loop;
end process;

----------------------------------------------------------------------------


end architecture behav;

