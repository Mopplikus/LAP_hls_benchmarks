    .INIT_00(256'h0250000504001f0102080d2055d2ff000206bc3240501f000250000401028000),
    .INIT_01(256'h0207b82056601001025000030bf2003302080d2055d280000207b2224072df02),
    .INIT_02(256'h02080d190012df020207c20b01f01f000250002f03b3207702080d0b00e20572),
    .INIT_03(256'h0207d00b0022202a001100202bb2202a001020202b22202a0250003641a28000),
    .INIT_04(256'h00bc0c0b0022202a00bd0d202c42202a00be0e324172202a00bf0f1d0022202a),
    .INIT_05(256'h001080207782202a020801202cd2202a025000324172202a0207fe1d0032202a),
    .INIT_06(256'h001100010822202a0010002f01f2202a0207d0224482202a001101010022202a),
    .INIT_07(256'h02500032439280000207151d0022df020207fe2200a01f010207ee205882202a),
    .INIT_08(256'h001101324391d0040010801d010320770207b2324391d0010208041d00820560),
    .INIT_09(256'h0207ee05040205630011002055d323ad0010043642b1d0080207d01d020322d6),
    .INIT_0A(256'h0208071d04020566025000224480106002072101002322d60207fe205661d004),
    .INIT_0B(256'h0207d02056620534001101030bf2052c0010802055d205720207b8364320109f),
    .INIT_0C(256'h0207fe3602a200370207ee1d08022bfc00110022448204fe0010080100220544),
    .INIT_0D(256'h0207c2010020900202080a2056625000025000030bf200630207322055d2004a),
    .INIT_0E(256'h00100c0b0020d0010207d02028c0b0000011012028332046001080224480d080),
    .INIT_0F(256'h0207470b0020121f0207fe20295011ff0207ee32443010ff0011001d00236046),
    .INIT_10(256'h036841207783e04000d0082029e1b20000900e324431b1000250001d00319001),
    .INIT_11(256'h032845010000d04000d002205660900100900e050402f0000250002055d01001),
    .INIT_12(256'h0328490900d2b00c00d0022200a2b00000900f205a0250000250002057232046),
    .INIT_13(256'h03284d0900d2d01000d00225000010ff0090103644b2bfff0250000d0802bf7e),
    .INIT_14(256'h032851014002d00100d002250000300f0090113644f090010250000d0402d011),
    .INIT_15(256'h00100c0b014090060008400b21536059000950013000d0200250000150b0900d),
    .INIT_16(256'h0131000d0080900d014808143000900601490e14200090060011000d01022054),
    .INIT_17(256'h036863011012205b01d10003007090070368591430036060019001142000d080),
    .INIT_18(256'h00d508224602054202500014106250000018ff3a464090070019ff1900109007),
    .INIT_19(256'h0018ff2d209205460019ff2d30a2050200110212350205360368691024020526),
    .INIT_1A(256'h00015001a002051e03e876250002054001d10302010205440250000900820534),
    .INIT_1B(256'h01410e09c1c2050201180114b06205080018ff14b06205480000400bb1320502),
    .INIT_1C(256'h00190b10ba00101901180809f1f2500003e86e09e1e204fe01400809d1d20506),
    .INIT_1D(256'h00084013f002022b00095013e002500002500013d003e07400110410cb019001),
    .INIT_1E(256'h0011022044b0d00103e87f204950900d01b90501b002021901981801a0420233),
    .INIT_1F(256'h0001802044b0108002500009d07206c30018ff2044b206bc0019ff09c073207a),
    .INIT_20(256'h01410601a731dc9301490009f07207fb0141062044b207d000381f09e0701101),
    .INIT_21(256'h0011020b612207e70149000b511010000141060b4100110001490001b013607d),
    .INIT_22(256'h01400612e601d11201400612d500311e000a9010c40001e0000080036012089c),
    .INIT_23(256'h0140063e4891d116014a001bb00320a401400619a011d11401400613f0032094),
    .INIT_24(256'h01d90b204952202a03d00001b01320c001da5d01a741d11a014a0025000320b2),
    .INIT_25(256'h0011042044f001e003a8992df07000d001d8142044f2f2390368972500001220),
    .INIT_26(256'h0250002044f1d05803a8972dd07030f801d8082044f140080250002de071410a),
    .INIT_27(256'h0095082044f1d08802f5032db07320ca0095082044f1d0480208b02dc07320ca),
    .INIT_28(256'h009508015002202a02f6050146c320cd02f504250001d0b80096082da07320cd),
    .INIT_29(256'h0095080d010001e002f6310b014000d002f5300b2152f2390096080130001220),
    .INIT_2A(256'h009508142001d04802f6380d008030f802f5371430014008009608142001410a),
    .INIT_2B(256'h025000190011d0b802f60601101320d002f53c030071d08800960814300320cd),
    .INIT_2C(256'h02d509102402f239001100224af01230001607141062202a0015ef3a4b3320d0),
    .INIT_2D(256'h00130009008140080250002d2091410a02d10b2d30a001e002d60a12350000d0),
    .INIT_2E(256'h02f0162d0081d0c80208d42d209320ca00b1172d30a1d08800b01606010030f8),
    .INIT_2F(256'h00b01814c002202a00130114b00320cd02f22014a061d0e802f11725000320cd),
    .INIT_30(256'h02f11925000001e002f01814f00000d00208d414e002f23900b11914d0001220),
    .INIT_31(256'h00b11b14c081d00800b01a14d08030f800130214e081400802f22114f0e1410a),
    .INIT_32(256'h02f222110b92f00202f11b250000100202f01a14a082202a0208d414b08320d0),
    .INIT_33(256'h0208d419011220d200b11d390002f00200b01c190e90100300130339000220d2),
    .INIT_34(256'h025000190f60120302f223390002021502f11d110072f00202f01c3e4d501004),
    .INIT_35(256'h03100000c000100101f1ff250002f03a01d0ff1100a01000001200250002f201),
    .INIT_36(256'h014006204df202590140062055220250014006204e920225014006204df2f024),
    .INIT_37(256'h01400e01100207fb01410025000202780140062055220247014100204e92023e),
    .INIT_38(256'h00b224141002027801003014c06207e701400e141000101001400e14c0601100),
    .INIT_39(256'h022bfc1410001100022bfc14c0620262022bfc141000110002500014c0601010),
    .INIT_3A(256'h022bfc11107206bc022bfc3a4ec207a4022bfc1d10a207e7022bfc2500001010),
    .INIT_3B(256'h022bfc2055501101022bfc01a0001080022bfc25000206bc022bfc1113020772),
    .INIT_3C(256'h022bfc0110401004022bfc3900001100022bfc204cb207fb022bfc09006207d0),
    .INIT_3D(256'h022bfc04a00207b2022bfc364f42023e022bfc19101207b2022bfc204bd207e7),
    .INIT_3E(256'h022bfc19201207b2022bfc2055220250022bfc204e9207b2022bfc0010020247),
    .INIT_3F(256'h022bfc22552206bc022bfc0110d20772022bfc25000206bc022bfc364ef20259),
    .INIT_40(256'h022bfc2255201014022bfc0115f01100022bfc22552207fb022bfc0112020278),
    .INIT_41(256'h022bfc22552207d0022bfc0113101101022bfc22552010c0022bfc0113e207e7),
    .INIT_42(256'h022bfc2255220262022bfc0113001100022bfc2255201014022bfc01133207b2),
    .INIT_43(256'h022bfc225520b002022bfc01132207e7022bfc2255201014022bfc0113101100),
    .INIT_44(256'h022bfc22552206bc022bfc01134207a4022bfc225523216b022bfc011331d002),
    .INIT_45(256'h022bfc22552206bc022bfc0113620772022bfc22552206bc022bfc0113520772),
    .INIT_46(256'h022bfc22552207fb022bfc01138207d0022bfc2255201101022bfc0113701080),
    .INIT_47(256'h022bfc22552207b8022bfc01141207e7022bfc2255201008022bfc0113901100),
    .INIT_48(256'h022bfc22552207b8022bfc0114320247022bfc22552207b8022bfc011422023e),
    .INIT_49(256'h022bfc22552206bc022bfc0114520259022bfc22552207b8022bfc0114420250),
    .INIT_4A(256'h022bfc22552206bc022bfc0114720772022bfc22552206bc022bfc0114620772),
    .INIT_4B(256'h022bfc2255201018022bfc0114901100022bfc22552207fb022bfc0114820278),
    .INIT_4C(256'h022bfc22552207d0022bfc0114b01101022bfc22552010c0022bfc0114a207e7),
    .INIT_4D(256'h022bfc2255220262022bfc0114d01100022bfc2255201018022bfc0114c207b8),
    .INIT_4E(256'h022bfc225520b002022bfc0114f207e7022bfc2255201018022bfc0114e01100),
    .INIT_4F(256'h022bfc22552206bc022bfc01151207a4022bfc225523216b022bfc011501d003),
    .INIT_50(256'h022bfc22552206bc022bfc0115320772022bfc22552206bc022bfc0115220772),
    .INIT_51(256'h022bfc2255201101022bfc0115501080022bfc22552206bc022bfc0115420772),
    .INIT_52(256'h022bfc225520100c022bfc0115701100022bfc22552207fb022bfc01156207d0),
    .INIT_53(256'h022bfc22552207c2022bfc011592023e022bfc22552207c2022bfc01158207e7),
    .INIT_54(256'h022bfc2d106207c2022bfc2055920250022bfc22552207c2022bfc0115a20247),
    .INIT_55(256'h022bfc36555206bc022bfc0d02020772022bfc0900d206bc022bfc2500020259),
    .INIT_56(256'h022bfc36559206bc022bfc0d01020772022bfc0900d206bc022bfc2500020772),
    .INIT_57(256'h022bfc250000101c022bfc0306001100022bfc09000207fb022bfc2500020278),
    .INIT_58(256'h022bfc09013207d0022bfc2500001101022bfc0309f010c0022bfc09000207e7),
    .INIT_59(256'h022bfc0316020262022bfc0010001100022bfc250000101c022bfc03007207c2),
    .INIT_5A(256'h022bfc20528206c9022bfc2d100207e7022bfc041000101c022bfc2056001100),
    .INIT_5B(256'h022bfc204d7207b2022bfc2055d206c9022bfc20500207b2022bfc20522206c6),
    .INIT_5C(256'h022bfc0319f3217f022bfc001001d002022bfc250000b002022bfc204fe206c6),
    .INIT_5D(256'h022bfc20542206c6022bfc2d100207b8022bfc04100206c9022bfc2055d207b8),
    .INIT_5E(256'h022bfc1d001207c2022bfc0b0323217f022bfc205001d003022bfc205220b002),
    .INIT_5F(256'h022bfc204fe202b2022bfc204d7206c6022bfc20560207c2022bfc3259c206c9),
    .INIT_60(256'h022bfc2050032189022bfc205221d002022bfc205420b002022bfc25000202bb),
    .INIT_61(256'h022bfc2500032189022bfc204fe1d003022bfc204d70b002022bfc01002202c4),
    .INIT_62(256'h022bfc0410001002022bfc2055d2b02e022bfc0319f20778022bfc00100202cd),
    .INIT_63(256'h022bfc2058801002022bfc010002d010022bfc2500001002022bfc2d1002d00f),
    .INIT_64(256'h022bfc2052220849022bfc205422b02e022bfc2d10320845022bfc0b1322d011),
    .INIT_65(256'h022bfc3259c1d002022bfc1d0010b002022bfc0b0322d00f022bfc2050001002),
    .INIT_66(256'h022bfc250002d010022bfc204fe01002022bfc204d72084d022bfc01040321a2),
    .INIT_67(256'h022bfc2500020851022bfc204fe321a2022bfc204d71d003022bfc010200b002),
    .INIT_68(256'h022bfc2053a2b02e022bfc325a720845022bfc1d0002d011022bfc2056001002),
    .INIT_69(256'h022bfc2052e0b002022bfc250002d00f022bfc2050001002022bfc2050420849),
    .INIT_6A(256'h022bfc2050001002022bfc205382084d022bfc20542321b3022bfc225a41d002),
    .INIT_6B(256'h022bfc20577321b3022bfc204fe1d003022bfc204d80b002022bfc00c302d010),
    .INIT_6C(256'h022bfc20500207a4022bfc2052e2d011022bfc2054001002022bfc2056b20851),
    .INIT_6D(256'h022bfc2500020278022bfc204fe206bc022bfc204d82021f022bfc0bc3a20215),
    .INIT_6E(256'h022bfc2050a01100022bfc205002026d022bfc2052801100022bfc2053601010),
    .INIT_6F(256'h022bfc0bc0520278022bfc204d8207b2022bfc0bc06207e7022bfc2050a01010),
    .INIT_70(256'h022bfc204fe01100022bfc204d82026d022bfc0bc0401100022bfc204d801014),
    .INIT_71(256'h022bfc205001d002022bfc205200b002022bfc20544207e7022bfc2060e01014),
    .INIT_72(256'h022bfc2062001018022bfc3a5cd20278022bfc0d504207b8022bfc09502321dc),
    .INIT_73(256'h022bfc09e1e01018022bfc09d1d01100022bfc09c1c2026d022bfc225e401100),
    .INIT_74(256'h022bfc14b06321dc022bfc14b061d003022bfc0bb130b002022bfc09f1f207e7),
    .INIT_75(256'h022bfc13f0001100022bfc13e000101c022bfc13d0020278022bfc10cb0207c2),
    .INIT_76(256'h022bfc2fc34207e7022bfc2fd350101c022bfc2fe3601100022bfc2ff3b2026d),
    .INIT_77(256'h022bfc204d80300f022bfc0bc3609001022bfc204d82b04e022bfc0bc3b20215),
    .INIT_78(256'h022bfc204d80d002022bfc0bc3409002022bfc204d832203022bfc0bc351d001),
    .INIT_79(256'h022bfc205002b40f022bfc205202b20f022bfc2052220778022bfc204fe321f4),
    .INIT_7A(256'h022bfc226022b10f022bfc206202b08f022bfc3a5ec2b04f022bfc0d5042b80f),
    .INIT_7B(256'h022bfc0bf3b2d010022bfc0be360101c022bfc0bd352d010022bfc0bc34010e0),
    .INIT_7C(256'h022bfc2044b2200a022bfc20495205a0022bfc01b0020572022bfc01a0401002),
    .INIT_7D(256'h022bfc2044b1d002022bfc09e070b002022bfc2044b2028c022bfc09f0720283),
    .INIT_7E(256'h022bfc204d81d003022bfc09c070b002022bfc2044b20295022bfc09d07321fe),
    .INIT_7F(256'h022bfc204d801000022bfc00ce020778022bfc204d82029e022bfc00cd0321fe),
    .INITP_00(256'h4952ce6a1e09d69332c842428bbab431f537b3fe77f060f076795bd6e453f1f2),
    .INITP_01(256'h406e489616f8128ffa7bfbd04b4d09ad44119b5dec49c1d04e172846ac067c4c),
    .INITP_02(256'hc225dc2cb38b1eb61b1632ffd42c1f4cfabb35d344099fcc6c9f0e58f428135b),
    .INITP_03(256'h2b6035a5986307243d19dea4330a7f0e07a724be8c7481472f3712eb00701c95),
    .INITP_04(256'h9f7718cbefda227895c1095a184f353aad3dba321d1e8ea08b3a351fa80595b9),
    .INITP_05(256'h352fc1dae7c61496a1616a4fda8fbe00764753a4964a629d83c54b809470d536),
    .INITP_06(256'h2b819fb90896870c57a007bb7ec96e73570920ae43d965d88eb5b9777eccc194),
    .INITP_07(256'h71c6f5efc6dacc7ef56c4168c3dac7504074f577e569f3f671d471dab3a88ba8),
    .INITP_08(256'hfae6fc52f7c275c9715b71da71cd764b7847f4cff4d5f4da7c4c7cc6f46bf742),
    .INITP_09(256'h717576f778fc75eff46e75787c6a7cfa7572f7617161717b71f3fa6dfaf9fa6f),
    .INITP_0A(256'h77615c7befe3417b6e6241727ac670e070ed70ff7af6f76675ec717e71e371f9),
    .INITP_0B(256'h4dd4c2ce436066f0cd7750524fecfc4c57d47473f272df4440f377c4c8f16954),
    .INITP_0C(256'heac245e6e0c949555b4b737268d26ddd4de5fae7524c4b707add57ebf2614efa),
    .INITP_0D(256'hf9577878fc7f78787bc6d1fbfeeed3c0cedd57c0727649ec71ee72f06f4ececc),
    .INITP_0E(256'h406b4ae16752516cf0d65dddfbe8c54efd78c452e142624fe56b4e65415ceadb),
    .INITP_0F(256'hd444dece454d62607be96fc8fd6fd1617e51c06b58f55ee46ef0f543d0f6dc68),
