`ifndef _DDR5MC_BFM_MAIN_REGS_DEFINE_VH_
`define _DDR5MC_BFM_MAIN_REGS_DEFINE_VH_

// spyglass disable_block ConstName
/* Address and Field defines*/

/* PCSR_LOCK */
`define DDRMC5_MAIN_PCSR_LOCK_OFFSET 16'hc
`define DDRMC5_MAIN_PCSR_LOCK_FLD_STATE 0
`define DDRMC5_MAIN_PCSR_LOCK_FLD_STATE_WIDTH 1
`define DDRMC5_MAIN_PCSR_LOCK_FLD_RESERVED 31:1
`define DDRMC5_MAIN_PCSR_LOCK_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_PCSR_LOCK_WIDTH 1

/* DDRMC_ECO */
`define DDRMC5_MAIN_DDRMC_ECO_OFFSET 16'h10
`define DDRMC5_MAIN_DDRMC_ECO_FLD_VAL 31:0
`define DDRMC5_MAIN_DDRMC_ECO_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_DDRMC_ECO_WIDTH 32

/* DDRMC_ISR */
`define DDRMC5_MAIN_DDRMC_ISR_OFFSET 16'h14
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_FATAL0 0
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_FATAL0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_FATAL1 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_FATAL1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CRYPTO_FATAL 2
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CRYPTO_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CRYPTO 3
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_0 4
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_1 5
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NSU_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_IN_LINE_ECC_0 6
`define DDRMC5_MAIN_DDRMC_ISR_FLD_IN_LINE_ECC_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_IN_LINE_ECC_1 7
`define DDRMC5_MAIN_DDRMC_ISR_FLD_IN_LINE_ECC_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_XMPU 8
`define DDRMC5_MAIN_DDRMC_ISR_FLD_XMPU_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CH0_DATA_PAR 9
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CH0_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CH1_DATA_PAR 10
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CH1_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC0_ECC0 11
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC1_ECC0 12
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC0_ECC1 13
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC1_ECC1 14
`define DDRMC5_MAIN_DDRMC_ISR_FLD_UC1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE0_ECC0 15
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE1_ECC0 16
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE0_ECC1 17
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE1_ECC1 18
`define DDRMC5_MAIN_DDRMC_ISR_FLD_CE1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD_FATAL 19
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD 20
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DC_CMD0_FATAL 21
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DC_CMD0_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_ADEC_PARITY_FATAL 22
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_ADEC_PARITY_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DC_CMD1_FATAL 23
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DC_CMD1_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD1 24
`define DDRMC5_MAIN_DDRMC_ISR_FLD_NA_CMD1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DRAM_PARITY0 25
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DRAM_PARITY0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_INTERNAL_PARITY 26
`define DDRMC5_MAIN_DDRMC_ISR_FLD_INTERNAL_PARITY_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DRAM_PARITY_FATAL_0 27
`define DDRMC5_MAIN_DDRMC_ISR_FLD_DRAM_PARITY_FATAL_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_SCAN_CLEAR_FAIL_CRYPTO 28
`define DDRMC5_MAIN_DDRMC_ISR_FLD_SCAN_CLEAR_FAIL_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_USER_0 29
`define DDRMC5_MAIN_DDRMC_ISR_FLD_USER_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_USER_1 30
`define DDRMC5_MAIN_DDRMC_ISR_FLD_USER_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_FLD_SCAN_CLEAR_FAIL 31
`define DDRMC5_MAIN_DDRMC_ISR_FLD_SCAN_CLEAR_FAIL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_ISR_WIDTH 32

/* DDRMC_ITR */
`define DDRMC5_MAIN_DDRMC_ITR_OFFSET 16'h18
`define DDRMC5_MAIN_DDRMC_ITR_WIDTH 32

/* DDRMC_IMR0 */
`define DDRMC5_MAIN_DDRMC_IMR0_OFFSET 16'h1c
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_FATAL0 0
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_FATAL0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_FATAL1 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_FATAL1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CRYPTO_FATAL 2
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CRYPTO_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CRYPTO 3
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_0 4
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_1 5
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NSU_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_IN_LINE_ECC_0 6
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_IN_LINE_ECC_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_IN_LINE_ECC_1 7
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_IN_LINE_ECC_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_XMPU 8
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_XMPU_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CH0_DATA_PAR 9
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CH0_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CH1_DATA_PAR 10
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CH1_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC0_ECC0 11
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC1_ECC0 12
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC0_ECC1 13
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC1_ECC1 14
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_UC1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE0_ECC0 15
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE1_ECC0 16
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE0_ECC1 17
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE1_ECC1 18
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_CE1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD_FATAL 19
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD 20
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DC_CMD0_FATAL 21
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DC_CMD0_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_ADEC_PARITY_FATAL 22
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_ADEC_PARITY_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DC_CMD1_FATAL 23
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DC_CMD1_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD1 24
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_NA_CMD1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DRAM_PARITY0 25
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DRAM_PARITY0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_INTERNAL_PARITY 26
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_INTERNAL_PARITY_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DRAM_PARITY_FATAL_0 27
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_DRAM_PARITY_FATAL_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_SCAN_CLEAR_FAIL_CRYPTO 28
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_SCAN_CLEAR_FAIL_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_USER_0 29
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_USER_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_USER_1 30
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_USER_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_SCAN_CLEAR_FAIL 31
`define DDRMC5_MAIN_DDRMC_IMR0_FLD_SCAN_CLEAR_FAIL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR0_WIDTH 32

/* DDRMC_IER0 */
`define DDRMC5_MAIN_DDRMC_IER0_OFFSET 16'h20
`define DDRMC5_MAIN_DDRMC_IER0_WIDTH 32

/* DDRMC_IDR0 */
`define DDRMC5_MAIN_DDRMC_IDR0_OFFSET 16'h24
`define DDRMC5_MAIN_DDRMC_IDR0_WIDTH 32

/* DDRMC_IMR1 */
`define DDRMC5_MAIN_DDRMC_IMR1_OFFSET 16'h28
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_FATAL0 0
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_FATAL0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_FATAL1 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_FATAL1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CRYPTO_FATAL 2
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CRYPTO_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CRYPTO 3
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_0 4
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_1 5
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NSU_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_IN_LINE_ECC_0 6
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_IN_LINE_ECC_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_IN_LINE_ECC_1 7
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_IN_LINE_ECC_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_XMPU 8
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_XMPU_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CH0_DATA_PAR 9
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CH0_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CH1_DATA_PAR 10
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CH1_DATA_PAR_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC0_ECC0 11
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC1_ECC0 12
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC0_ECC1 13
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC1_ECC1 14
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_UC1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE0_ECC0 15
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE0_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE1_ECC0 16
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE1_ECC0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE0_ECC1 17
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE0_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE1_ECC1 18
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_CE1_ECC1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD_FATAL 19
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD 20
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DC_CMD0_FATAL 21
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DC_CMD0_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_ADEC_PARITY_FATAL 22
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_ADEC_PARITY_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DC_CMD1_FATAL 23
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DC_CMD1_FATAL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD1 24
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_NA_CMD1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DRAM_PARITY0 25
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DRAM_PARITY0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_INTERNAL_PARITY 26
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_INTERNAL_PARITY_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DRAM_PARITY_FATAL_0 27
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_DRAM_PARITY_FATAL_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_SCAN_CLEAR_FAIL_CRYPTO 28
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_SCAN_CLEAR_FAIL_CRYPTO_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_USER_0 29
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_USER_0_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_USER_1 30
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_USER_1_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_SCAN_CLEAR_FAIL 31
`define DDRMC5_MAIN_DDRMC_IMR1_FLD_SCAN_CLEAR_FAIL_WIDTH 1
`define DDRMC5_MAIN_DDRMC_IMR1_WIDTH 32

/* DDRMC_IER1 */
`define DDRMC5_MAIN_DDRMC_IER1_OFFSET 16'h2c
`define DDRMC5_MAIN_DDRMC_IER1_WIDTH 32

/* DDRMC_IDR1 */
`define DDRMC5_MAIN_DDRMC_IDR1_OFFSET 16'h30
`define DDRMC5_MAIN_DDRMC_IDR1_WIDTH 32

/* DDRMC_IOR */
`define DDRMC5_MAIN_DDRMC_IOR_OFFSET 16'h34
`define DDRMC5_MAIN_DDRMC_IOR_FLD_OFFSET 4:0
`define DDRMC5_MAIN_DDRMC_IOR_FLD_OFFSET_WIDTH 5
`define DDRMC5_MAIN_DDRMC_IOR_FLD_RESERVED 31:5
`define DDRMC5_MAIN_DDRMC_IOR_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_DDRMC_IOR_WIDTH 5

/* REG_REF_3 */
`define DDRMC5_MAIN_REG_REF_3_OFFSET 16'h200
`define DDRMC5_MAIN_REG_REF_3_FLD_AFTER_ZQ_WAIT_TIME 9:0
`define DDRMC5_MAIN_REG_REF_3_FLD_AFTER_ZQ_WAIT_TIME_WIDTH 10
`define DDRMC5_MAIN_REG_REF_3_FLD_BEFORE_ZQ_WAIT_TIME 19:10
`define DDRMC5_MAIN_REG_REF_3_FLD_BEFORE_ZQ_WAIT_TIME_WIDTH 10
`define DDRMC5_MAIN_REG_REF_3_FLD_RESERVED 31:20
`define DDRMC5_MAIN_REG_REF_3_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_REG_REF_3_WIDTH 20

/* REG_REF_4 */
`define DDRMC5_MAIN_REG_REF_4_OFFSET 16'h204
`define DDRMC5_MAIN_REG_REF_4_FLD_LPDDR4_REFRESH_TYPE 0
`define DDRMC5_MAIN_REG_REF_4_FLD_LPDDR4_REFRESH_TYPE_WIDTH 1
`define DDRMC5_MAIN_REG_REF_4_FLD_REFRESH_FORCE_IN_RR 1
`define DDRMC5_MAIN_REG_REF_4_FLD_REFRESH_FORCE_IN_RR_WIDTH 1
`define DDRMC5_MAIN_REG_REF_4_FLD_RESERVED 31:2
`define DDRMC5_MAIN_REG_REF_4_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_REG_REF_4_WIDTH 2

/* REG_REF_5 */
`define DDRMC5_MAIN_REG_REF_5_OFFSET 16'h208
`define DDRMC5_MAIN_REG_REF_5_FLD_DDR5_ECS_ENABLE 0
`define DDRMC5_MAIN_REG_REF_5_FLD_DDR5_ECS_ENABLE_WIDTH 1
`define DDRMC5_MAIN_REG_REF_5_FLD_TREFI_BASED_ECS_TIMER 20:1
`define DDRMC5_MAIN_REG_REF_5_FLD_TREFI_BASED_ECS_TIMER_WIDTH 20
`define DDRMC5_MAIN_REG_REF_5_FLD_RESERVED 31:21
`define DDRMC5_MAIN_REG_REF_5_FLD_RESERVED_WIDTH 11
`define DDRMC5_MAIN_REG_REF_5_WIDTH 21

/* REG_SCRUB_TO */
`define DDRMC5_MAIN_REG_SCRUB_TO_OFFSET 16'h20c
`define DDRMC5_MAIN_REG_SCRUB_TO_FLD_SCRUB_TIMEOUT_INTVL 31:0
`define DDRMC5_MAIN_REG_SCRUB_TO_FLD_SCRUB_TIMEOUT_INTVL_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_TO_WIDTH 32

/* REG_TXN_CONFIG */
`define DDRMC5_MAIN_REG_TXN_CONFIG_OFFSET 16'h210
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_STARVED_TIMER 15:0
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_STARVED_TIMER_WIDTH 16
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_ALL_CMD_ARB_MODE 16
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_ALL_CMD_ARB_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_ARB_ONLY_MODE 17
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_ARB_ONLY_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_AND_STARVED_ARB_ONLY_MODE 18
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_AND_STARVED_ARB_ONLY_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_WR_PRI_ARB_ONLY_MODE 19
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_TXNQ_RD_PRI_WR_PRI_ARB_ONLY_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PH_BLOCK_EN 20
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PH_BLOCK_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_CMD_PRI_BUS_DIR_EN 21
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_CMD_PRI_BUS_DIR_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PM_BLOCK_EN 22
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PM_BLOCK_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PC_BLOCK_EN 23
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_PC_BLOCK_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_AGE_BLOCK_EN 24
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_AGE_BLOCK_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_WAR_MODE 26:25
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_WAR_MODE_WIDTH 2
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_RESERVED 31:27
`define DDRMC5_MAIN_REG_TXN_CONFIG_FLD_RESERVED_WIDTH 5
`define DDRMC5_MAIN_REG_TXN_CONFIG_WIDTH 27

/* REG_TXN_CONFIG_1 */
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_OFFSET 16'h214
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_TXNQ_SKIP_FRAC_EN 0
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_TXNQ_SKIP_FRAC_EN_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_TXNQ_OTHER_CAS_COMPARE_WR_ONLY 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_TXNQ_OTHER_CAS_COMPARE_WR_ONLY_WIDTH 1
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_HI_INC 5:2
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_HI_INC_WIDTH 4
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_MID_INC 9:6
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_MID_INC_WIDTH 4
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_LOW_INC 13:10
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_LOW_INC_WIDTH 4
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_DEFAULT_INC 17:14
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_DEFAULT_INC_WIDTH 4
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_HI_THRESHOLD 24:18
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_HI_THRESHOLD_WIDTH 7
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_MID_THRESHOLD 31:25
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_FLD_SKIP_MID_THRESHOLD_WIDTH 7
`define DDRMC5_MAIN_REG_TXN_CONFIG_1_WIDTH 32

/* REG_TXN_CONFIG_2 */
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_OFFSET 16'h218
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_FLD_SKIP_LOW_THRESHOLD 6:0
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_FLD_SKIP_LOW_THRESHOLD_WIDTH 7
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_FLD_RESERVED 31:7
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_REG_TXN_CONFIG_2_WIDTH 7

/* REG_TXN_CONFIG_3 */
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_OFFSET 16'h21c
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_FLD_TXNQ_STARVED_MODE_TIMER 15:0
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_FLD_TXNQ_STARVED_MODE_TIMER_WIDTH 16
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_TXN_CONFIG_3_WIDTH 16

/* REG_WR_CONFIG */
`define DDRMC5_MAIN_REG_WR_CONFIG_OFFSET 16'h220
`define DDRMC5_MAIN_REG_WR_CONFIG_FLD_TXNQ_WR_RD_PRI_TIMER 15:0
`define DDRMC5_MAIN_REG_WR_CONFIG_FLD_TXNQ_WR_RD_PRI_TIMER_WIDTH 16
`define DDRMC5_MAIN_REG_WR_CONFIG_FLD_TXNQ_WR_TOP_TIMER 31:16
`define DDRMC5_MAIN_REG_WR_CONFIG_FLD_TXNQ_WR_TOP_TIMER_WIDTH 16
`define DDRMC5_MAIN_REG_WR_CONFIG_WIDTH 32

/* REG_RD_CONFIG */
`define DDRMC5_MAIN_REG_RD_CONFIG_OFFSET 16'h224
`define DDRMC5_MAIN_REG_RD_CONFIG_FLD_FULL_THRESHOLD 5:0
`define DDRMC5_MAIN_REG_RD_CONFIG_FLD_FULL_THRESHOLD_WIDTH 6
`define DDRMC5_MAIN_REG_RD_CONFIG_FLD_RESERVED 31:6
`define DDRMC5_MAIN_REG_RD_CONFIG_FLD_RESERVED_WIDTH 26
`define DDRMC5_MAIN_REG_RD_CONFIG_WIDTH 6

/* REG_PT_CONFIG */
`define DDRMC5_MAIN_REG_PT_CONFIG_OFFSET 16'h228
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PAGE_POLICY 1:0
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PAGE_POLICY_WIDTH 2
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PT_BGRL_MODE 3:2
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PT_BGRL_MODE_WIDTH 2
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PAGE_TIMER 19:4
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_PAGE_TIMER_WIDTH 16
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_RESERVED 31:20
`define DDRMC5_MAIN_REG_PT_CONFIG_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_REG_PT_CONFIG_WIDTH 20

/* REG_DRAM_ARB */
`define DDRMC5_MAIN_REG_DRAM_ARB_OFFSET 16'h22c
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_WRITE_LEVEL_HI 4:0
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_WRITE_LEVEL_HI_WIDTH 5
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_RESERVED 7:5
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_RESERVED_WIDTH 3
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_WRITE_LEVEL_LO 12:8
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_WRITE_LEVEL_LO_WIDTH 5
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_RESERVED_1 31:13
`define DDRMC5_MAIN_REG_DRAM_ARB_FLD_RESERVED_1_WIDTH 19
`define DDRMC5_MAIN_REG_DRAM_ARB_WIDTH 13

/* REG_CONFIG0 */
`define DDRMC5_MAIN_REG_CONFIG0_OFFSET 16'h230
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DRAM_TYPE 0
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DRAM_TYPE_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DDR4_2T 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DDR4_2T_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DDR5_SDR_ADDR 2
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DDR5_SDR_ADDR_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED 3
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DRAM_WIDTH 5:4
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DRAM_WIDTH_WIDTH 2
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED_1 11:6
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DIMM_TYPE 13:12
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DIMM_TYPE_WIDTH 2
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_RANKS 15:14
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_RANKS_WIDTH 2
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_SLOTS 16
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_SLOTS_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_CH 17
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_CH_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_WIDTH_PER_CH 19:18
`define DDRMC5_MAIN_REG_CONFIG0_FLD_WIDTH_PER_CH_WIDTH 2
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_LRANKS 22:20
`define DDRMC5_MAIN_REG_CONFIG0_FLD_NUM_LRANKS_WIDTH 3
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DM_EN 23
`define DDRMC5_MAIN_REG_CONFIG0_FLD_DM_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_BYPASS_AFTER_PARTIAL_WR_EN 24
`define DDRMC5_MAIN_REG_CONFIG0_FLD_BYPASS_AFTER_PARTIAL_WR_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_AUTO_PRECHARGE_EN 25
`define DDRMC5_MAIN_REG_CONFIG0_FLD_AUTO_PRECHARGE_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_SPLIT_ACT_EN 26
`define DDRMC5_MAIN_REG_CONFIG0_FLD_SPLIT_ACT_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_PH_BLOCK_EN 27
`define DDRMC5_MAIN_REG_CONFIG0_FLD_PH_BLOCK_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_CMD_PRI_BUS_DIR_EN 28
`define DDRMC5_MAIN_REG_CONFIG0_FLD_CMD_PRI_BUS_DIR_EN_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED_2 31:29
`define DDRMC5_MAIN_REG_CONFIG0_FLD_RESERVED_2_WIDTH 3
`define DDRMC5_MAIN_REG_CONFIG0_WIDTH 29

/* REG_PINOUT */
`define DDRMC5_MAIN_REG_PINOUT_OFFSET 16'h234
`define DDRMC5_MAIN_REG_PINOUT_FLD_PO_SELECT 4:0
`define DDRMC5_MAIN_REG_PINOUT_FLD_PO_SELECT_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_ENCODE_EN 5
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_ENCODE_EN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_CORRECT_EN 6
`define DDRMC5_MAIN_REG_PINOUT_FLD_CORRECT_EN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_IO_ENABLE 7
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_IO_ENABLE_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED 9:8
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_POISON_BIT_EN 10
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_POISON_BIT_EN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_ADDR_PAR_EN 11
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_ADDR_PAR_EN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_BURST_ORDER_EN 12
`define DDRMC5_MAIN_REG_PINOUT_FLD_ECC_BURST_ORDER_EN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED_1 13
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_DIMM_CHAN 14
`define DDRMC5_MAIN_REG_PINOUT_FLD_DIMM_CHAN_WIDTH 1
`define DDRMC5_MAIN_REG_PINOUT_FLD_SWAP_CK 18:15
`define DDRMC5_MAIN_REG_PINOUT_FLD_SWAP_CK_WIDTH 4
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED_2 31:19
`define DDRMC5_MAIN_REG_PINOUT_FLD_RESERVED_2_WIDTH 13
`define DDRMC5_MAIN_REG_PINOUT_WIDTH 19

/* REG_PINOUT_ADDR_MUX_0 */
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_OFFSET 16'h238
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR0 4:0
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR0_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR1 9:5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR1_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR2 14:10
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR2_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR3 19:15
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR3_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR4 24:20
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR4_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR5 29:25
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_ADDR5_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_0_WIDTH 30

/* REG_PINOUT_ADDR_MUX_1 */
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_OFFSET 16'h23c
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR6 4:0
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR6_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR7 9:5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR7_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR8 14:10
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR8_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR9 19:15
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR9_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR10 24:20
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR10_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR11 29:25
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_ADDR11_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_1_WIDTH 30

/* REG_PINOUT_ADDR_MUX_2 */
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_OFFSET 16'h240
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_ADDR12 4:0
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_ADDR12_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_ADDR13 9:5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_ADDR13_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS0 14:10
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS0_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS1 19:15
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS1_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS2 24:20
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS2_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS3 29:25
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_CS3_WIDTH 5
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_PINOUT_ADDR_MUX_2_WIDTH 30

/* REG_CONFIG3 */
`define DDRMC5_MAIN_REG_CONFIG3_OFFSET 16'h244
`define DDRMC5_MAIN_REG_CONFIG3_FLD_SPARE 15:0
`define DDRMC5_MAIN_REG_CONFIG3_FLD_SPARE_WIDTH 16
`define DDRMC5_MAIN_REG_CONFIG3_FLD_SPARE2 31:16
`define DDRMC5_MAIN_REG_CONFIG3_FLD_SPARE2_WIDTH 16
`define DDRMC5_MAIN_REG_CONFIG3_WIDTH 32

/* REG_CONFIG4 */
`define DDRMC5_MAIN_REG_CONFIG4_OFFSET 16'h248
`define DDRMC5_MAIN_REG_CONFIG4_FLD_SPARE 19:0
`define DDRMC5_MAIN_REG_CONFIG4_FLD_SPARE_WIDTH 20
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RROB_RETURN_DLY 22:20
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RROB_RETURN_DLY_WIDTH 3
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RROB_RETURN_MODE 23
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RROB_RETURN_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RESERVED 31:24
`define DDRMC5_MAIN_REG_CONFIG4_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_REG_CONFIG4_WIDTH 24

/* A2A_DUAL_CHAN */
`define DDRMC5_MAIN_A2A_DUAL_CHAN_OFFSET 16'h24c
`define DDRMC5_MAIN_A2A_DUAL_CHAN_FLD_EN 0
`define DDRMC5_MAIN_A2A_DUAL_CHAN_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_A2A_DUAL_CHAN_FLD_RESERVED 31:1
`define DDRMC5_MAIN_A2A_DUAL_CHAN_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_A2A_DUAL_CHAN_WIDTH 1

/* A2A_RD_MAP */
`define DDRMC5_MAIN_A2A_RD_MAP_OFFSET 16'h250
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_ALERT 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_ALERT_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_LBDQ 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_LBDQ_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_RESERVED 31:14
`define DDRMC5_MAIN_A2A_RD_MAP_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_A2A_RD_MAP_WIDTH 14

/* A2A_RD_MAP_DQ_0 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_OFFSET 16'h254
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL0 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL0_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL1 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL1_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL2 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL2_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL3 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_MUX_CNTRL3_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_0_WIDTH 28

/* A2A_RD_MAP_DQ_1 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_OFFSET 16'h258
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL4 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL4_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL5 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL5_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL6 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL6_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL7 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_MUX_CNTRL7_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_1_WIDTH 28

/* A2A_RD_MAP_DQ_2 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_OFFSET 16'h25c
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL8 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL8_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL9 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL9_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL10 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL10_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL11 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_MUX_CNTRL11_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_2_WIDTH 28

/* A2A_RD_MAP_DQ_3 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_OFFSET 16'h260
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL12 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL12_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL13 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL13_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL14 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL14_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL15 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_MUX_CNTRL15_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_3_WIDTH 28

/* A2A_RD_MAP_DQ_4 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_OFFSET 16'h264
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL16 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL16_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL17 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL17_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL18 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL18_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL19 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_MUX_CNTRL19_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_4_WIDTH 28

/* A2A_RD_MAP_DQ_5 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_OFFSET 16'h268
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL20 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL20_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL21 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL21_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL22 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL22_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL23 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_MUX_CNTRL23_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_5_WIDTH 28

/* A2A_RD_MAP_DQ_6 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_OFFSET 16'h26c
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL24 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL24_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL25 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL25_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL26 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL26_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL27 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_MUX_CNTRL27_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_6_WIDTH 28

/* A2A_RD_MAP_DQ_7 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_OFFSET 16'h270
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL28 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL28_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL29 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL29_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL30 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL30_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL31 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_MUX_CNTRL31_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_7_WIDTH 28

/* A2A_RD_MAP_DQ_8 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_OFFSET 16'h274
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL32 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL32_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL33 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL33_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL34 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL34_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL35 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_MUX_CNTRL35_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_8_WIDTH 28

/* A2A_RD_MAP_DQ_9 */
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_OFFSET 16'h278
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL36 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL36_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL37 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL37_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL38 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL38_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL39 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_MUX_CNTRL39_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DQ_9_WIDTH 28

/* A2A_RD_MAP_DBI_CH0_0 */
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_OFFSET 16'h27c
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL0 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL0_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL1 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL1_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL2 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL2_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL3 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_MUX_CNTRL3_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_0_WIDTH 28

/* A2A_RD_MAP_DBI_CH0_1 */
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_OFFSET 16'h280
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_FLD_MUX_CNTRL4 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_FLD_MUX_CNTRL4_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_FLD_RESERVED 31:7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH0_1_WIDTH 7

/* A2A_RD_MAP_DBI_CH1_0 */
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_OFFSET 16'h284
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL0 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL0_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL1 13:7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL1_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL2 20:14
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL2_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL3 27:21
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_MUX_CNTRL3_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_0_WIDTH 28

/* A2A_RD_MAP_DBI_CH1_1 */
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_OFFSET 16'h288
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_FLD_MUX_CNTRL4 6:0
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_FLD_MUX_CNTRL4_WIDTH 7
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_RD_MAP_DBI_CH1_1_WIDTH 7

/* A2A_PIN_MAP_0 */
`define DDRMC5_MAIN_A2A_PIN_MAP_0_OFFSET 16'h28c
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL0 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL0_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL1 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL1_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL2 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL2_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL3 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_MUX_CNTRL3_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_0_WIDTH 28

/* A2A_PIN_MAP_1 */
`define DDRMC5_MAIN_A2A_PIN_MAP_1_OFFSET 16'h290
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL4 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL4_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL5 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL5_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL6 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL6_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL7 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_MUX_CNTRL7_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_1_WIDTH 28

/* A2A_PIN_MAP_2 */
`define DDRMC5_MAIN_A2A_PIN_MAP_2_OFFSET 16'h294
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL8 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL8_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL9 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL9_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL10 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL10_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL11 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_MUX_CNTRL11_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_2_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_2_WIDTH 28

/* A2A_PIN_MAP_3 */
`define DDRMC5_MAIN_A2A_PIN_MAP_3_OFFSET 16'h298
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL12 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL12_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL13 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL13_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL14 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL14_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL15 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_MUX_CNTRL15_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_3_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_3_WIDTH 28

/* A2A_PIN_MAP_4 */
`define DDRMC5_MAIN_A2A_PIN_MAP_4_OFFSET 16'h29c
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL16 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL16_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL17 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL17_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL18 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL18_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL19 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_MUX_CNTRL19_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_4_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_4_WIDTH 28

/* A2A_PIN_MAP_5 */
`define DDRMC5_MAIN_A2A_PIN_MAP_5_OFFSET 16'h2a0
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL20 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL20_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL21 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL21_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL22 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL22_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL23 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_MUX_CNTRL23_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_5_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_5_WIDTH 28

/* A2A_PIN_MAP_6 */
`define DDRMC5_MAIN_A2A_PIN_MAP_6_OFFSET 16'h2a4
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL24 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL24_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL25 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL25_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL26 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL26_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL27 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_MUX_CNTRL27_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_6_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_6_WIDTH 28

/* A2A_PIN_MAP_7 */
`define DDRMC5_MAIN_A2A_PIN_MAP_7_OFFSET 16'h2a8
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL28 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL28_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL29 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL29_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL30 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL30_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL31 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_MUX_CNTRL31_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_7_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_7_WIDTH 28

/* A2A_PIN_MAP_8 */
`define DDRMC5_MAIN_A2A_PIN_MAP_8_OFFSET 16'h2ac
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL32 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL32_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL33 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL33_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL34 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL34_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL35 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_MUX_CNTRL35_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_8_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_8_WIDTH 28

/* A2A_PIN_MAP_9 */
`define DDRMC5_MAIN_A2A_PIN_MAP_9_OFFSET 16'h2b0
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL36 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL36_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL37 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL37_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL38 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL38_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL39 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_MUX_CNTRL39_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_9_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_9_WIDTH 28

/* A2A_PIN_MAP_10 */
`define DDRMC5_MAIN_A2A_PIN_MAP_10_OFFSET 16'h2b4
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL40 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL40_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL41 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL41_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL42 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL42_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL43 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_MUX_CNTRL43_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_10_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_10_WIDTH 28

/* A2A_PIN_MAP_11 */
`define DDRMC5_MAIN_A2A_PIN_MAP_11_OFFSET 16'h2b8
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL44 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL44_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL45 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL45_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL46 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL46_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL47 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_MUX_CNTRL47_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_11_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_11_WIDTH 28

/* A2A_PIN_MAP_12 */
`define DDRMC5_MAIN_A2A_PIN_MAP_12_OFFSET 16'h2bc
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL48 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL48_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL49 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL49_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL50 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL50_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL51 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_MUX_CNTRL51_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_12_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_12_WIDTH 28

/* A2A_PIN_MAP_13 */
`define DDRMC5_MAIN_A2A_PIN_MAP_13_OFFSET 16'h2c0
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL52 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL52_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL53 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL53_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL54 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL54_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL55 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_MUX_CNTRL55_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_13_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_13_WIDTH 28

/* A2A_PIN_MAP_14 */
`define DDRMC5_MAIN_A2A_PIN_MAP_14_OFFSET 16'h2c4
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL56 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL56_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL57 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL57_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL58 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL58_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL59 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_MUX_CNTRL59_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_14_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_14_WIDTH 28

/* A2A_PIN_MAP_15 */
`define DDRMC5_MAIN_A2A_PIN_MAP_15_OFFSET 16'h2c8
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL60 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL60_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL61 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL61_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL62 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL62_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL63 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_MUX_CNTRL63_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_15_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_15_WIDTH 28

/* A2A_PIN_MAP_16 */
`define DDRMC5_MAIN_A2A_PIN_MAP_16_OFFSET 16'h2cc
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL64 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL64_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL65 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL65_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL66 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL66_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL67 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_MUX_CNTRL67_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_16_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_16_WIDTH 28

/* A2A_PIN_MAP_17 */
`define DDRMC5_MAIN_A2A_PIN_MAP_17_OFFSET 16'h2d0
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL68 6:0
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL68_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL69 13:7
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL69_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL70 20:14
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL70_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL71 27:21
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_MUX_CNTRL71_WIDTH 7
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_RESERVED 31:28
`define DDRMC5_MAIN_A2A_PIN_MAP_17_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_A2A_PIN_MAP_17_WIDTH 28

/* A2A_DIFF_T_PIN_MAP_0 */
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_OFFSET 16'h2d4
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL0 5:0
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL0_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL1 11:6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL1_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL2 17:12
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL2_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL3 23:18
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL3_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL4 29:24
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_MUX_CNTRL4_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_0_WIDTH 30

/* A2A_DIFF_T_PIN_MAP_1 */
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_OFFSET 16'h2d8
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL5 5:0
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL5_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL6 11:6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL6_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL7 17:12
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL7_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL8 23:18
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL8_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL9 29:24
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_MUX_CNTRL9_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_1_WIDTH 30

/* A2A_DIFF_T_PIN_MAP_2 */
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_OFFSET 16'h2dc
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_MUX_CNTRL10 5:0
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_MUX_CNTRL10_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_MUX_CNTRL11 11:6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_MUX_CNTRL11_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_RESERVED 31:12
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_A2A_DIFF_T_PIN_MAP_2_WIDTH 12

/* A2A_DIFF_C_PIN_MAP_0 */
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_OFFSET 16'h2e0
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL0 5:0
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL0_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL1 11:6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL1_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL2 17:12
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL2_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL3 23:18
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL3_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL4 29:24
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_MUX_CNTRL4_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_0_WIDTH 30

/* A2A_DIFF_C_PIN_MAP_1 */
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_OFFSET 16'h2e4
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL5 5:0
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL5_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL6 11:6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL6_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL7 17:12
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL7_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL8 23:18
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL8_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL9 29:24
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_MUX_CNTRL9_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_1_WIDTH 30

/* A2A_DIFF_C_PIN_MAP_2 */
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_OFFSET 16'h2e8
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_MUX_CNTRL10 5:0
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_MUX_CNTRL10_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_MUX_CNTRL11 11:6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_MUX_CNTRL11_WIDTH 6
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_RESERVED 31:12
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_A2A_DIFF_C_PIN_MAP_2_WIDTH 12

/* A2A_CNTRL_MAP_0 */
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_OFFSET 16'h2ec
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL0 5:0
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL0_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL1 11:6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL1_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL2 17:12
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL2_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL3 23:18
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL3_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL4 29:24
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_MUX_CNTRL4_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_CNTRL_MAP_0_WIDTH 30

/* A2A_CNTRL_MAP_1 */
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_OFFSET 16'h2f0
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL5 5:0
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL5_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL6 11:6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL6_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL7 17:12
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL7_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL8 23:18
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL8_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL9 29:24
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_MUX_CNTRL9_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_A2A_CNTRL_MAP_1_WIDTH 30

/* A2A_CNTRL_MAP_2 */
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_OFFSET 16'h2f4
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_MUX_CNTRL10 5:0
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_MUX_CNTRL10_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_MUX_CNTRL11 11:6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_MUX_CNTRL11_WIDTH 6
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_RESERVED 31:12
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_A2A_CNTRL_MAP_2_WIDTH 12

/* XPI_MAP_PD_EN */
`define DDRMC5_MAIN_XPI_MAP_PD_EN_OFFSET 16'h2f8
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB0 3:0
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB0_WIDTH 4
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB1 7:4
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB1_WIDTH 4
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB2 11:8
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_HB2_WIDTH 4
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_RESERVED 31:12
`define DDRMC5_MAIN_XPI_MAP_PD_EN_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_XPI_MAP_PD_EN_WIDTH 12

/* RAM_SETTING_RF2PHS */
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_OFFSET 16'h2fc
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMAA 2:0
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMAA_WIDTH 3
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMAB 5:3
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMAB_WIDTH 3
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMASA 6
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_EMASA_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_STOV 7
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_STOV_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_RESERVED 31:8
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_RAM_SETTING_RF2PHS_WIDTH 8

/* RAM_SETTING_SRSPHD */
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_OFFSET 16'h300
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMA 2:0
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMA_WIDTH 3
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMAW 4:3
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMAW_WIDTH 2
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMAS 5
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_EMAS_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_STOV 6
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_STOV_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_RESERVED 31:7
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_RAM_SETTING_SRSPHD_WIDTH 7

/* RAM_SETTING_RFSPHD */
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_OFFSET 16'h304
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMA 2:0
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMA_WIDTH 3
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMAW 4:3
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMAW_WIDTH 2
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMAS 5
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_EMAS_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_STOV 6
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_STOV_WIDTH 1
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_RESERVED 31:7
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_RAM_SETTING_RFSPHD_WIDTH 7

/* LP5_MRS_BIT_MUX_BYTE0 */
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_OFFSET 16'h308
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT0 2:0
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT0_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT1 5:3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT1_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT2 8:6
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT2_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT3 11:9
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT3_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT4 14:12
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT4_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT5 17:15
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT5_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT6 20:18
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT6_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT7 23:21
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_BIT7_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_RESERVED 31:24
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE0_WIDTH 24

/* LP5_MRS_BIT_MUX_BYTE1 */
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_OFFSET 16'h30c
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT0 2:0
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT0_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT1 5:3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT1_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT2 8:6
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT2_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT3 11:9
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT3_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT4 14:12
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT4_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT5 17:15
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT5_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT6 20:18
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT6_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT7 23:21
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_BIT7_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_RESERVED 31:24
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE1_WIDTH 24

/* LP5_MRS_BIT_MUX_BYTE2 */
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_OFFSET 16'h310
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT0 2:0
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT0_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT1 5:3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT1_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT2 8:6
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT2_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT3 11:9
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT3_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT4 14:12
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT4_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT5 17:15
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT5_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT6 20:18
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT6_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT7 23:21
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_BIT7_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_RESERVED 31:24
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE2_WIDTH 24

/* LP5_MRS_BIT_MUX_BYTE3 */
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_OFFSET 16'h314
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT0 2:0
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT0_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT1 5:3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT1_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT2 8:6
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT2_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT3 11:9
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT3_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT4 14:12
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT4_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT5 17:15
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT5_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT6 20:18
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT6_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT7 23:21
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_BIT7_WIDTH 3
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_RESERVED 31:24
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_LP5_MRS_BIT_MUX_BYTE3_WIDTH 24

/* TXNQ_RD_PRIORITY */
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_OFFSET 16'h318
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_LOW 7:0
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_LOW_WIDTH 8
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_MED 15:8
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_MED_WIDTH 8
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_HIGH 23:16
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_TH_HIGH_WIDTH 8
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_SKIP_COUNT_EN 24
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_SKIP_COUNT_EN_WIDTH 1
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_ONLY_READ 25
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_ONLY_READ_WIDTH 1
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_RESERVED 31:26
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_FLD_RESERVED_WIDTH 6
`define DDRMC5_MAIN_TXNQ_RD_PRIORITY_WIDTH 26

/* TXNQ_WR_PRIORITY */
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_OFFSET 16'h31c
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_LOW 7:0
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_LOW_WIDTH 8
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_MED 15:8
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_MED_WIDTH 8
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_HIGH 23:16
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_TH_HIGH_WIDTH 8
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_SKIP_COUNT_EN 24
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_SKIP_COUNT_EN_WIDTH 1
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_RESERVED 31:25
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_FLD_RESERVED_WIDTH 7
`define DDRMC5_MAIN_TXNQ_WR_PRIORITY_WIDTH 25

/* TXNQ_ENTRY_COUNT_MODE */
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_OFFSET 16'h320
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_ENABLE 0
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_ENABLE_WIDTH 1
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_RESERVED 3:1
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_RESERVED_WIDTH 3
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_LIMIT 13:4
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_LIMIT_WIDTH 10
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_RESERVED_1 31:14
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_FLD_RESERVED_1_WIDTH 18
`define DDRMC5_MAIN_TXNQ_ENTRY_COUNT_MODE_WIDTH 14

/* DDR5_SPARE_STA_CFG0 */
`define DDRMC5_MAIN_DDR5_SPARE_STA_CFG0_OFFSET 16'h324
`define DDRMC5_MAIN_DDR5_SPARE_STA_CFG0_FLD_SPARE 31:0
`define DDRMC5_MAIN_DDR5_SPARE_STA_CFG0_FLD_SPARE_WIDTH 32
`define DDRMC5_MAIN_DDR5_SPARE_STA_CFG0_WIDTH 32

/* REG_SAFE_CONFIG0 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_OFFSET 16'h800
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TCCD_S_SR 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TCCD_S_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TCCD_L_SR 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TCCD_L_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TRRD_S 20:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TRRD_S_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TRRD_L 25:21
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_TRRD_L_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_RESERVED 31:26
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_FLD_RESERVED_WIDTH 6
`define DDRMC5_MAIN_REG_SAFE_CONFIG0_WIDTH 26

/* REG_SAFE_CONFIG1 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_OFFSET 16'h804
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_R2R_DR 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_R2R_DR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_R2R_SR_DLR 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_R2R_SR_DLR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_W2W_DR 23:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_W2W_DR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_W2W_SR_DLR 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_FLD_TCS_W2W_SR_DLR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG1_WIDTH 32

/* REG_SAFE_CONFIG2 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_OFFSET 16'h808
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRCD 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRCD_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRP 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRP_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRAS 23:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TRAS_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TFAW_DLR 29:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_TFAW_DLR_WIDTH 6
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_SAFE_CONFIG2_WIDTH 30

/* REG_SAFE_CONFIG3 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_OFFSET 16'h80c
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_L_SR 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_L_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_S_SR 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_S_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_DR 23:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_DR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_SR_DLR 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_FLD_TCS_W2R_SR_DLR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG3_WIDTH 32

/* REG_SAFE_CONFIG4 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_OFFSET 16'h810
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TRTP 4:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TRTP_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_R2W_SR 12:5
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_R2W_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_R2W_DR 20:13
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_R2W_DR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_W2P 28:21
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_TCS_W2P_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_RESERVED 31:29
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_FLD_RESERVED_WIDTH 3
`define DDRMC5_MAIN_REG_SAFE_CONFIG4_WIDTH 29

/* REG_SAFE_CONFIG5 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_OFFSET 16'h814
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_CAS_LATENCY 6:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_CAS_LATENCY_WIDTH 7
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_RESERVED 7
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_CWL 14:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_CWL_WIDTH 7
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_TRP_AB 22:15
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_TRP_AB_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_RESERVED_1 27:23
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_RESERVED_1_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_ADD_CMD_DELAY 30:28
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_ADD_CMD_DELAY_WIDTH 3
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_ADD_CMD_DELAY_EN 31
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_FLD_ADD_CMD_DELAY_EN_WIDTH 1
`define DDRMC5_MAIN_REG_SAFE_CONFIG5_WIDTH 32

/* REG_SAFE_CONFIG6 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_OFFSET 16'h818
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TREFI 15:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TREFI_WIDTH 16
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TPBR2PBR 25:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TPBR2PBR_WIDTH 10
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TPBR2ACT 30:26
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_TPBR2ACT_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_RESERVED 31
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_REG_SAFE_CONFIG6_WIDTH 31

/* REG_SAFE_CONFIG7 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_OFFSET 16'h81c
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_SLR_AB 11:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_SLR_AB_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_DLR_PB 23:12
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_DLR_PB_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_R2R 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_FLD_TRFC_R2R_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG7_WIDTH 32

/* REG_SAFE_CONFIG8 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG8_OFFSET 16'h820
`define DDRMC5_MAIN_REG_SAFE_CONFIG8_FLD_TZQCS_ITVL_REFI_BASED 31:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG8_FLD_TZQCS_ITVL_REFI_BASED_WIDTH 32
`define DDRMC5_MAIN_REG_SAFE_CONFIG8_WIDTH 32

/* REG_SAFE_CONFIG9 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_OFFSET 16'h824
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCD_L_WR 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCD_L_WR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCD_L_WR2 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCD_L_WR2_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCS_R2W_S_SR 23:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCS_R2W_S_SR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCDMW 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_FLD_TCCDMW_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG9_WIDTH 32

/* REG_SAFE_CONFIG10 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_OFFSET 16'h828
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TIMING_DERATE_CYCLES 4:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TIMING_DERATE_CYCLES_WIDTH 5
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_RESERVED 19:5
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TRRD_DLR 23:20
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TRRD_DLR_WIDTH 4
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TFAW 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_FLD_TFAW_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG10_WIDTH 32

/* REG_SAFE_CONFIG11 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_OFFSET 16'h82c
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TREFSBRD_SLR 7:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TREFSBRD_SLR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TREFSBRD_DLR 15:8
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TREFSBRD_DLR_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TRFC_DPR 27:16
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_TRFC_DPR_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_RESERVED 31:28
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_REG_SAFE_CONFIG11_WIDTH 28

/* REG_SAFE_CONFIG12 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_OFFSET 16'h830
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_TRFM_AB 11:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_TRFM_AB_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_TRFM_PB 23:12
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_TRFM_PB_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_RESERVED 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG12_WIDTH 24

/* REG_SAFE_CONFIG13 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_OFFSET 16'h834
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_TRFC_SB_SLR 11:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_TRFC_SB_SLR_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_TRFC_SB_DLR 23:12
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_TRFC_SB_DLR_WIDTH 12
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_RESERVED 31:24
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_REG_SAFE_CONFIG13_WIDTH 24

/* REG_SAFE_CONFIG14 */
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_OFFSET 16'h838
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RDA2ACT_SB 9:0
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RDA2ACT_SB_WIDTH 10
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RESERVED 11:10
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_WRA2ACT_SB 21:12
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_WRA2ACT_SB_WIDTH 10
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RESERVED_1 31:22
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_FLD_RESERVED_1_WIDTH 10
`define DDRMC5_MAIN_REG_SAFE_CONFIG14_WIDTH 22

/* REG_SAFE_MUX */
`define DDRMC5_MAIN_REG_SAFE_MUX_OFFSET 16'h83c
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_SELECT 0
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_SELECT_WIDTH 1
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_TIMING_DERATE_EN 1
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_TIMING_DERATE_EN_WIDTH 1
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_RESERVED 31:2
`define DDRMC5_MAIN_REG_SAFE_MUX_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_REG_SAFE_MUX_WIDTH 2

/* REG_RETRY_0 */
`define DDRMC5_MAIN_REG_RETRY_0_OFFSET 16'h840
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE 2:0
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE_WIDTH 3
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE2 7:3
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE2_WIDTH 5
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE3 15:8
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE3_WIDTH 8
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE4 22:16
`define DDRMC5_MAIN_REG_RETRY_0_FLD_SPARE4_WIDTH 7
`define DDRMC5_MAIN_REG_RETRY_0_FLD_RMW_FIFO_DEALLOC_PERIOD 28:23
`define DDRMC5_MAIN_REG_RETRY_0_FLD_RMW_FIFO_DEALLOC_PERIOD_WIDTH 6
`define DDRMC5_MAIN_REG_RETRY_0_FLD_RESERVED 31:29
`define DDRMC5_MAIN_REG_RETRY_0_FLD_RESERVED_WIDTH 3
`define DDRMC5_MAIN_REG_RETRY_0_WIDTH 29

/* REG_RETRY_1 */
`define DDRMC5_MAIN_REG_RETRY_1_OFFSET 16'h844
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RETRY_WAIT_TIMER 6:0
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RETRY_WAIT_TIMER_WIDTH 7
`define DDRMC5_MAIN_REG_RETRY_1_FLD_REF_EXTRA_NUM 9:7
`define DDRMC5_MAIN_REG_RETRY_1_FLD_REF_EXTRA_NUM_WIDTH 3
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE 10
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE_WIDTH 1
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE2 16:11
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE2_WIDTH 6
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE3 17
`define DDRMC5_MAIN_REG_RETRY_1_FLD_SPARE3_WIDTH 1
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RETRY_FIFO_DEALLOC_PERIOD 23:18
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RETRY_FIFO_DEALLOC_PERIOD_WIDTH 6
`define DDRMC5_MAIN_REG_RETRY_1_FLD_WR_FIFO_DEALLOC_PERIOD 29:24
`define DDRMC5_MAIN_REG_RETRY_1_FLD_WR_FIFO_DEALLOC_PERIOD_WIDTH 6
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_REG_RETRY_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_RETRY_1_WIDTH 30

/* REG_RETRY_2 */
`define DDRMC5_MAIN_REG_RETRY_2_OFFSET 16'h848
`define DDRMC5_MAIN_REG_RETRY_2_FLD_READ_FIFO_DEALLOC_PERIOD 5:0
`define DDRMC5_MAIN_REG_RETRY_2_FLD_READ_FIFO_DEALLOC_PERIOD_WIDTH 6
`define DDRMC5_MAIN_REG_RETRY_2_FLD_RESERVED 7:6
`define DDRMC5_MAIN_REG_RETRY_2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_RETRY_2_FLD_HS_WATCHDOG 27:8
`define DDRMC5_MAIN_REG_RETRY_2_FLD_HS_WATCHDOG_WIDTH 20
`define DDRMC5_MAIN_REG_RETRY_2_FLD_HS_WATCHDOG_EN 28
`define DDRMC5_MAIN_REG_RETRY_2_FLD_HS_WATCHDOG_EN_WIDTH 1
`define DDRMC5_MAIN_REG_RETRY_2_FLD_RESERVED_1 31:29
`define DDRMC5_MAIN_REG_RETRY_2_FLD_RESERVED_1_WIDTH 3
`define DDRMC5_MAIN_REG_RETRY_2_WIDTH 29

/* REG_REF_0 */
`define DDRMC5_MAIN_REG_REF_0_OFFSET 16'h84c
`define DDRMC5_MAIN_REG_REF_0_FLD_REFRESH_SPEED 2:0
`define DDRMC5_MAIN_REG_REF_0_FLD_REFRESH_SPEED_WIDTH 3
`define DDRMC5_MAIN_REG_REF_0_FLD_RESERVED 31:3
`define DDRMC5_MAIN_REG_REF_0_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_REG_REF_0_WIDTH 3

/* REG_REF_1 */
`define DDRMC5_MAIN_REG_REF_1_OFFSET 16'h850
`define DDRMC5_MAIN_REG_REF_1_FLD_TZQLAT 7:0
`define DDRMC5_MAIN_REG_REF_1_FLD_TZQLAT_WIDTH 8
`define DDRMC5_MAIN_REG_REF_1_FLD_TZQ_START_LATCH_ITVL 20:8
`define DDRMC5_MAIN_REG_REF_1_FLD_TZQ_START_LATCH_ITVL_WIDTH 13
`define DDRMC5_MAIN_REG_REF_1_FLD_RESERVED 31:21
`define DDRMC5_MAIN_REG_REF_1_FLD_RESERVED_WIDTH 11
`define DDRMC5_MAIN_REG_REF_1_WIDTH 21

/* REG_REF_2 */
`define DDRMC5_MAIN_REG_REF_2_OFFSET 16'h854
`define DDRMC5_MAIN_REG_REF_2_FLD_TRAFFIC_BASED_SELFREFRESH_EN 0
`define DDRMC5_MAIN_REG_REF_2_FLD_TRAFFIC_BASED_SELFREFRESH_EN_WIDTH 1
`define DDRMC5_MAIN_REG_REF_2_FLD_TRAFFIC_BASED_POWERDOWN_EN 1
`define DDRMC5_MAIN_REG_REF_2_FLD_TRAFFIC_BASED_POWERDOWN_EN_WIDTH 1
`define DDRMC5_MAIN_REG_REF_2_FLD_PDE_ODT_EN 2
`define DDRMC5_MAIN_REG_REF_2_FLD_PDE_ODT_EN_WIDTH 1
`define DDRMC5_MAIN_REG_REF_2_FLD_RESERVED 31:3
`define DDRMC5_MAIN_REG_REF_2_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_REG_REF_2_WIDTH 3

/* REG_COM_1 */
`define DDRMC5_MAIN_REG_COM_1_OFFSET 16'h858
`define DDRMC5_MAIN_REG_COM_1_FLD_T_IDLE_ITVL_SELFREFRESH 26:0
`define DDRMC5_MAIN_REG_COM_1_FLD_T_IDLE_ITVL_SELFREFRESH_WIDTH 27
`define DDRMC5_MAIN_REG_COM_1_FLD_RESERVED 31:27
`define DDRMC5_MAIN_REG_COM_1_FLD_RESERVED_WIDTH 5
`define DDRMC5_MAIN_REG_COM_1_WIDTH 27

/* REG_COM_2 */
`define DDRMC5_MAIN_REG_COM_2_OFFSET 16'h85c
`define DDRMC5_MAIN_REG_COM_2_FLD_T_IDLE_ITVL_POWERDOWN 26:0
`define DDRMC5_MAIN_REG_COM_2_FLD_T_IDLE_ITVL_POWERDOWN_WIDTH 27
`define DDRMC5_MAIN_REG_COM_2_FLD_RESERVED 31:27
`define DDRMC5_MAIN_REG_COM_2_FLD_RESERVED_WIDTH 5
`define DDRMC5_MAIN_REG_COM_2_WIDTH 27

/* REG_COM_3 */
`define DDRMC5_MAIN_REG_COM_3_OFFSET 16'h860
`define DDRMC5_MAIN_REG_COM_3_FLD_TCSPD 5:0
`define DDRMC5_MAIN_REG_COM_3_FLD_TCSPD_WIDTH 6
`define DDRMC5_MAIN_REG_COM_3_FLD_TXP 11:6
`define DDRMC5_MAIN_REG_COM_3_FLD_TXP_WIDTH 6
`define DDRMC5_MAIN_REG_COM_3_FLD_TCACSH 14:12
`define DDRMC5_MAIN_REG_COM_3_FLD_TCACSH_WIDTH 3
`define DDRMC5_MAIN_REG_COM_3_FLD_TCSH 17:15
`define DDRMC5_MAIN_REG_COM_3_FLD_TCSH_WIDTH 3
`define DDRMC5_MAIN_REG_COM_3_FLD_T_BLOCK_DRAIN_OUT 23:18
`define DDRMC5_MAIN_REG_COM_3_FLD_T_BLOCK_DRAIN_OUT_WIDTH 6
`define DDRMC5_MAIN_REG_COM_3_FLD_T_SR_ENTRY_WAIT 31:24
`define DDRMC5_MAIN_REG_COM_3_FLD_T_SR_ENTRY_WAIT_WIDTH 8
`define DDRMC5_MAIN_REG_COM_3_WIDTH 32

/* REG_MRS_0 */
`define DDRMC5_MAIN_REG_MRS_0_OFFSET 16'h864
`define DDRMC5_MAIN_REG_MRS_0_FLD_TCS_MRW_2_ANY 5:0
`define DDRMC5_MAIN_REG_MRS_0_FLD_TCS_MRW_2_ANY_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_0_FLD_TCS_MRR_2_ANY 11:6
`define DDRMC5_MAIN_REG_MRS_0_FLD_TCS_MRR_2_ANY_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_0_FLD_TOSCI_START_2_READ 25:12
`define DDRMC5_MAIN_REG_MRS_0_FLD_TOSCI_START_2_READ_WIDTH 14
`define DDRMC5_MAIN_REG_MRS_0_FLD_RESERVED 31:26
`define DDRMC5_MAIN_REG_MRS_0_FLD_RESERVED_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_0_WIDTH 26

/* REG_MRS_1 */
`define DDRMC5_MAIN_REG_MRS_1_OFFSET 16'h868
`define DDRMC5_MAIN_REG_MRS_1_FLD_TOSCI_CMD_ITVL 25:0
`define DDRMC5_MAIN_REG_MRS_1_FLD_TOSCI_CMD_ITVL_WIDTH 26
`define DDRMC5_MAIN_REG_MRS_1_FLD_TCS_MPC_2_ANY 31:26
`define DDRMC5_MAIN_REG_MRS_1_FLD_TCS_MPC_2_ANY_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_1_WIDTH 32

/* REG_MRS_2 */
`define DDRMC5_MAIN_REG_MRS_2_OFFSET 16'h86c
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN 0
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN_LPDDR5_1 1
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN_LPDDR5_1_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_2_FLD_RESERVED 2
`define DDRMC5_MAIN_REG_MRS_2_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN_ALL_RANK 3
`define DDRMC5_MAIN_REG_MRS_2_FLD_MRS_OSCI_EN_ALL_RANK_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_2_FLD_RESERVED_1 31:4
`define DDRMC5_MAIN_REG_MRS_2_FLD_RESERVED_1_WIDTH 28
`define DDRMC5_MAIN_REG_MRS_2_WIDTH 4

/* REG_MRS_7 */
`define DDRMC5_MAIN_REG_MRS_7_OFFSET 16'h870
`define DDRMC5_MAIN_REG_MRS_7_FLD_T_MR_BLOCK_ITVL 11:0
`define DDRMC5_MAIN_REG_MRS_7_FLD_T_MR_BLOCK_ITVL_WIDTH 12
`define DDRMC5_MAIN_REG_MRS_7_FLD_RESERVED 31:12
`define DDRMC5_MAIN_REG_MRS_7_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_REG_MRS_7_WIDTH 12

/* REG_SCRUB_INTVL */
`define DDRMC5_MAIN_REG_SCRUB_INTVL_OFFSET 16'h874
`define DDRMC5_MAIN_REG_SCRUB_INTVL_FLD_SCRUB_INTVL 23:0
`define DDRMC5_MAIN_REG_SCRUB_INTVL_FLD_SCRUB_INTVL_WIDTH 24
`define DDRMC5_MAIN_REG_SCRUB_INTVL_FLD_RESERVED 31:24
`define DDRMC5_MAIN_REG_SCRUB_INTVL_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_REG_SCRUB_INTVL_WIDTH 24

/* REG_SCRUB_TAP */
`define DDRMC5_MAIN_REG_SCRUB_TAP_OFFSET 16'h878
`define DDRMC5_MAIN_REG_SCRUB_TAP_FLD_SCRUB_INTVL_TAP 23:0
`define DDRMC5_MAIN_REG_SCRUB_TAP_FLD_SCRUB_INTVL_TAP_WIDTH 24
`define DDRMC5_MAIN_REG_SCRUB_TAP_FLD_RESERVED 31:24
`define DDRMC5_MAIN_REG_SCRUB_TAP_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_REG_SCRUB_TAP_WIDTH 24

/* REG_SCRUB_PER_RD */
`define DDRMC5_MAIN_REG_SCRUB_PER_RD_OFFSET 16'h87c
`define DDRMC5_MAIN_REG_SCRUB_PER_RD_FLD_PERIODIC_READ_INTVL 31:0
`define DDRMC5_MAIN_REG_SCRUB_PER_RD_FLD_PERIODIC_READ_INTVL_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_PER_RD_WIDTH 32

/* REG_SCRUB_CONFIG */
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_OFFSET 16'h880
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_SCRUB_FILL_MODE 0
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_SCRUB_FILL_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_SCRUB_LOOP_MODE 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_SCRUB_LOOP_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_PERIODIC_READ_INTVL_EN 2
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_PERIODIC_READ_INTVL_EN_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_ON_DIE_EN 3
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_ON_DIE_EN_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_PER_RANK_NA_PER_RD 4
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_PER_RANK_NA_PER_RD_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_RESERVED 31:5
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_REG_SCRUB_CONFIG_WIDTH 5

/* REG_SCRUB_OTF */
`define DDRMC5_MAIN_REG_SCRUB_OTF_OFFSET 16'h884
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_OTF_SCRUB_EN_0 0
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_OTF_SCRUB_EN_0_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_OTF_SCRUB_EN_1 1
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_OTF_SCRUB_EN_1_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_RESERVED 31:2
`define DDRMC5_MAIN_REG_SCRUB_OTF_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_REG_SCRUB_OTF_WIDTH 2

/* REG_SCRUB_BASE_ADDR_LO */
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_LO_OFFSET 16'h888
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_LO_FLD_SCRUB_BASE_ADDR_ON_DIE 31:0
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_LO_FLD_SCRUB_BASE_ADDR_ON_DIE_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_LO_WIDTH 32

/* REG_SCRUB_BASE_ADDR_HI */
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_OFFSET 16'h88c
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_FLD_SCRUB_BASE_ADDR_ON_DIE 15:0
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_FLD_SCRUB_BASE_ADDR_ON_DIE_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_BASE_ADDR_HI_WIDTH 16

/* REG_SCRUB_ADDR_RANGE_LO */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_LO_OFFSET 16'h890
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_LO_FLD_SCRUB_ADDR_RANGE_ON_DIE 31:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_LO_FLD_SCRUB_ADDR_RANGE_ON_DIE_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_LO_WIDTH 32

/* REG_SCRUB_ADDR_RANGE_HI */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_OFFSET 16'h894
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_FLD_SCRUB_ADDR_RANGE_ON_DIE 3:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_FLD_SCRUB_ADDR_RANGE_ON_DIE_WIDTH 4
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_SCRUB_ADDR_RANGE_HI_WIDTH 4

/* REG_SCRUB_DEBUG_MODE */
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_OFFSET 16'h898
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_SCRUB_DEBUG_MODE_0 0
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_SCRUB_DEBUG_MODE_0_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_SCRUB_DEBUG_MODE_1 1
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_SCRUB_DEBUG_MODE_1_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_RESERVED 31:2
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_REG_SCRUB_DEBUG_MODE_WIDTH 2

/* REG_RFM */
`define DDRMC5_MAIN_REG_RFM_OFFSET 16'h89c
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_EN 0
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_EN_WIDTH 1
`define DDRMC5_MAIN_REG_RFM_FLD_RAAIMT 5:1
`define DDRMC5_MAIN_REG_RFM_FLD_RAAIMT_WIDTH 5
`define DDRMC5_MAIN_REG_RFM_FLD_RAAMULT 8:6
`define DDRMC5_MAIN_REG_RFM_FLD_RAAMULT_WIDTH 3
`define DDRMC5_MAIN_REG_RFM_FLD_RAADEC_REF 11:9
`define DDRMC5_MAIN_REG_RFM_FLD_RAADEC_REF_WIDTH 3
`define DDRMC5_MAIN_REG_RFM_FLD_RAADEC_RFM 14:12
`define DDRMC5_MAIN_REG_RFM_FLD_RAADEC_RFM_WIDTH 3
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_MODE 15
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_ACT_HOLD_TH 26:16
`define DDRMC5_MAIN_REG_RFM_FLD_RFM_ACT_HOLD_TH_WIDTH 11
`define DDRMC5_MAIN_REG_RFM_FLD_FGR_MODE 27
`define DDRMC5_MAIN_REG_RFM_FLD_FGR_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_RFM_FLD_RESERVED 31:28
`define DDRMC5_MAIN_REG_RFM_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_REG_RFM_WIDTH 28

/* REG_RFM_1 */
`define DDRMC5_MAIN_REG_RFM_1_OFFSET 16'h8a0
`define DDRMC5_MAIN_REG_RFM_1_FLD_RFM_TRIGGER_TH 10:0
`define DDRMC5_MAIN_REG_RFM_1_FLD_RFM_TRIGGER_TH_WIDTH 11
`define DDRMC5_MAIN_REG_RFM_1_FLD_RESERVED 31:11
`define DDRMC5_MAIN_REG_RFM_1_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_REG_RFM_1_WIDTH 11

/* REG_CONFIG1 */
`define DDRMC5_MAIN_REG_CONFIG1_OFFSET 16'h8a4
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_MODE 0
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_MODE_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_EN_0 1
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_EN_0_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_EN_1 2
`define DDRMC5_MAIN_REG_CONFIG1_FLD_REF_EN_1_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG1_FLD_RESERVED 31:3
`define DDRMC5_MAIN_REG_CONFIG1_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_REG_CONFIG1_WIDTH 3

/* REG_CONFIG2 */
`define DDRMC5_MAIN_REG_CONFIG2_OFFSET 16'h8a8
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED 0
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED_1 20:1
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED_1_WIDTH 20
`define DDRMC5_MAIN_REG_CONFIG2_FLD_PER_RD_H_THRESH 30:21
`define DDRMC5_MAIN_REG_CONFIG2_FLD_PER_RD_H_THRESH_WIDTH 10
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED_2 31
`define DDRMC5_MAIN_REG_CONFIG2_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_MAIN_REG_CONFIG2_WIDTH 31

/* CAL_MODE */
`define DDRMC5_MAIN_CAL_MODE_OFFSET 16'h8ac
`define DDRMC5_MAIN_CAL_MODE_FLD_BYPASS 0
`define DDRMC5_MAIN_CAL_MODE_FLD_BYPASS_WIDTH 1
`define DDRMC5_MAIN_CAL_MODE_FLD_RESERVED 31:1
`define DDRMC5_MAIN_CAL_MODE_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_CAL_MODE_WIDTH 1

/* X5PHYIO_STARTUP */
`define DDRMC5_MAIN_X5PHYIO_STARTUP_OFFSET 16'h8b0
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_RST 0
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_RST_WIDTH 1
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_WRCS 1
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_WRCS_WIDTH 1
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_CONFIG_RANK 3:2
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_CONFIG_RANK_WIDTH 2
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_CONFIG_SLOT 7:4
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_CONFIG_SLOT_WIDTH 4
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_RESERVED 31:8
`define DDRMC5_MAIN_X5PHYIO_STARTUP_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_X5PHYIO_STARTUP_WIDTH 8

/* XPI_DQS_T_CNTRL_PREAMBLE0 */
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE0_OFFSET 16'h8b4
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE0_FLD_PATTERN 31:0
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE0_FLD_PATTERN_WIDTH 32
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE0_WIDTH 32

/* XPI_DQS_T_CNTRL_PREAMBLE1 */
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE1_OFFSET 16'h8b8
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE1_FLD_PATTERN 31:0
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE1_FLD_PATTERN_WIDTH 32
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_PREAMBLE1_WIDTH 32

/* XPI_DQS_T_CNTRL */
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_OFFSET 16'h8bc
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_BURST_PATTERN 15:0
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_BURST_PATTERN_WIDTH 16
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_POSTAMBLE_PATTERN 23:16
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_POSTAMBLE_PATTERN_WIDTH 8
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_RESERVED 31:24
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_XPI_DQS_T_CNTRL_WIDTH 24

/* XPI_OE_CNTRL_PREAMBLE */
`define DDRMC5_MAIN_XPI_OE_CNTRL_PREAMBLE_OFFSET 16'h8c0
`define DDRMC5_MAIN_XPI_OE_CNTRL_PREAMBLE_FLD_PATTERN 31:0
`define DDRMC5_MAIN_XPI_OE_CNTRL_PREAMBLE_FLD_PATTERN_WIDTH 32
`define DDRMC5_MAIN_XPI_OE_CNTRL_PREAMBLE_WIDTH 32

/* XPI_OE_CNTRL */
`define DDRMC5_MAIN_XPI_OE_CNTRL_OFFSET 16'h8c4
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_BURST_PATTERN 7:0
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_BURST_PATTERN_WIDTH 8
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_POSTAMBLE_PATTERN 11:8
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_POSTAMBLE_PATTERN_WIDTH 4
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED 15:12
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_PREAMBLE_LENGTH_TCK 20:16
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_PREAMBLE_LENGTH_TCK_WIDTH 5
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_1 21
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_POSTAMBLE_LENGTH_TCK 24:22
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_POSTAMBLE_LENGTH_TCK_WIDTH 3
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_2 26:25
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_2_WIDTH 2
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RD_PREAMBLE_LENGTH_TCK 30:27
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RD_PREAMBLE_LENGTH_TCK_WIDTH 4
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_3 31
`define DDRMC5_MAIN_XPI_OE_CNTRL_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_MAIN_XPI_OE_CNTRL_WIDTH 31

/* XPI_OE_CNTRL2 */
`define DDRMC5_MAIN_XPI_OE_CNTRL2_OFFSET 16'h8c8
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_RESERVED 0
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_WRCS_EARLY 2:1
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_WRCS_EARLY_WIDTH 2
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_DQS_DQ_DM_1CLK_LATE 3
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_DQS_DQ_DM_1CLK_LATE_WIDTH 1
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_RESERVED_1 31:4
`define DDRMC5_MAIN_XPI_OE_CNTRL2_FLD_RESERVED_1_WIDTH 28
`define DDRMC5_MAIN_XPI_OE_CNTRL2_WIDTH 4

/* DBG_TRIGGER */
`define DDRMC5_MAIN_DBG_TRIGGER_OFFSET 16'h8cc
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_EN 0
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_SOURCE 2:1
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_SOURCE_WIDTH 2
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_RESERVED 31:3
`define DDRMC5_MAIN_DBG_TRIGGER_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_DBG_TRIGGER_WIDTH 3

/* CAL_CS_CH */
`define DDRMC5_MAIN_CAL_CS_CH_OFFSET 16'h8d0
`define DDRMC5_MAIN_CAL_CS_CH_FLD_EN 0
`define DDRMC5_MAIN_CAL_CS_CH_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_CAL_CS_CH_FLD_SEL 1
`define DDRMC5_MAIN_CAL_CS_CH_FLD_SEL_WIDTH 1
`define DDRMC5_MAIN_CAL_CS_CH_FLD_CS_NOP 2
`define DDRMC5_MAIN_CAL_CS_CH_FLD_CS_NOP_WIDTH 1
`define DDRMC5_MAIN_CAL_CS_CH_FLD_RESERVED 31:3
`define DDRMC5_MAIN_CAL_CS_CH_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_CAL_CS_CH_WIDTH 3

/* XPI_MAP_CS_OVERRIDE_CFG */
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_OFFSET 16'h8d4
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_CH0_EN 0
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_CH0_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_CH1_EN 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_CH1_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_RESERVED 31:2
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_CFG_WIDTH 2

/* XPI_OE_ALL_NIB */
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_OFFSET 16'h8d8
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_DLY 6:0
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_DLY_WIDTH 7
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_DLY_OFFSET 10:7
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_DLY_OFFSET_WIDTH 4
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_RESERVED 31:11
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_XPI_OE_ALL_NIB_WIDTH 11

/* XPI_WRDATA_ALL_NIB */
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_OFFSET 16'h8dc
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DLY 6:0
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DLY_WIDTH 7
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DLY_OFFSET 10:7
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DLY_OFFSET_WIDTH 4
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_SHIFT_180DEG 11
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_SHIFT_180DEG_WIDTH 1
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DQ_IDLE 12
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DQ_IDLE_WIDTH 1
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DM_IDLE 13
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DM_IDLE_WIDTH 1
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DQS_T_IDLE 14
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_DQS_T_IDLE_WIDTH 1
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_RESERVED 31:15
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_FLD_RESERVED_WIDTH 17
`define DDRMC5_MAIN_XPI_WRDATA_ALL_NIB_WIDTH 15

/* XPI_PMI_CONFIG */
`define DDRMC5_MAIN_XPI_PMI_CONFIG_OFFSET 16'h8e0
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_PAR_EN 0
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_PAR_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_ALERT_EN 1
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_ALERT_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_RESERVED 31:2
`define DDRMC5_MAIN_XPI_PMI_CONFIG_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_XPI_PMI_CONFIG_WIDTH 2

/* XPI_WRITE_DM_DBI */
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_OFFSET 16'h8e4
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_CFG_EN 1:0
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_CFG_EN_WIDTH 2
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_RESERVED 3:2
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_DM_INVERT 4
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_DM_INVERT_WIDTH 1
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_RESERVED_1 31:5
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_FLD_RESERVED_1_WIDTH 27
`define DDRMC5_MAIN_XPI_WRITE_DM_DBI_WIDTH 5

/* XPI_WRITE_NIB_ENABLE */
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_OFFSET 16'h8e8
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_FLD_SEL 9:0
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_FLD_SEL_WIDTH 10
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_XPI_WRITE_NIB_ENABLE_WIDTH 10

/* CK_PATTERN */
`define DDRMC5_MAIN_CK_PATTERN_OFFSET 16'h8ec
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_T 7:0
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_T_WIDTH 8
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_N 15:8
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_N_WIDTH 8
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_MODE 16
`define DDRMC5_MAIN_CK_PATTERN_FLD_CK_MODE_WIDTH 1
`define DDRMC5_MAIN_CK_PATTERN_FLD_RESERVED 31:17
`define DDRMC5_MAIN_CK_PATTERN_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_CK_PATTERN_WIDTH 17

/* PRBS_SEED0 */
`define DDRMC5_MAIN_PRBS_SEED0_OFFSET 16'h8f0
`define DDRMC5_MAIN_PRBS_SEED0_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED0_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED0_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED0_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED0_WIDTH 23

/* PRBS_SEED1 */
`define DDRMC5_MAIN_PRBS_SEED1_OFFSET 16'h8f4
`define DDRMC5_MAIN_PRBS_SEED1_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED1_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED1_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED1_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED1_WIDTH 23

/* PRBS_SEED2 */
`define DDRMC5_MAIN_PRBS_SEED2_OFFSET 16'h8f8
`define DDRMC5_MAIN_PRBS_SEED2_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED2_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED2_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED2_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED2_WIDTH 23

/* PRBS_SEED3 */
`define DDRMC5_MAIN_PRBS_SEED3_OFFSET 16'h8fc
`define DDRMC5_MAIN_PRBS_SEED3_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED3_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED3_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED3_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED3_WIDTH 23

/* PRBS_SEED4 */
`define DDRMC5_MAIN_PRBS_SEED4_OFFSET 16'h900
`define DDRMC5_MAIN_PRBS_SEED4_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED4_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED4_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED4_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED4_WIDTH 23

/* PRBS_SEED5 */
`define DDRMC5_MAIN_PRBS_SEED5_OFFSET 16'h904
`define DDRMC5_MAIN_PRBS_SEED5_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED5_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED5_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED5_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED5_WIDTH 23

/* PRBS_SEED6 */
`define DDRMC5_MAIN_PRBS_SEED6_OFFSET 16'h908
`define DDRMC5_MAIN_PRBS_SEED6_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED6_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED6_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED6_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED6_WIDTH 23

/* PRBS_SEED7 */
`define DDRMC5_MAIN_PRBS_SEED7_OFFSET 16'h90c
`define DDRMC5_MAIN_PRBS_SEED7_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED7_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED7_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED7_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED7_WIDTH 23

/* PRBS_SEED8 */
`define DDRMC5_MAIN_PRBS_SEED8_OFFSET 16'h910
`define DDRMC5_MAIN_PRBS_SEED8_FLD_DATA 22:0
`define DDRMC5_MAIN_PRBS_SEED8_FLD_DATA_WIDTH 23
`define DDRMC5_MAIN_PRBS_SEED8_FLD_RESERVED 31:23
`define DDRMC5_MAIN_PRBS_SEED8_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_PRBS_SEED8_WIDTH 23

/* PHY_RANK_WRITE_OVERRIDE */
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_OFFSET 16'h914
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_STATIC_ENABLE 1:0
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_STATIC_ENABLE_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK0 3:2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK0_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK1 5:4
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK1_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK2 7:6
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK2_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK3 9:8
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH0_RANK3_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK0 11:10
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK0_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK1 13:12
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK1_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK2 15:14
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK2_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK3 17:16
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_CH1_RANK3_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_RESERVED 31:18
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_WIDTH 18

/* CLK_GATE */
`define DDRMC5_MAIN_CLK_GATE_OFFSET 16'h918
`define DDRMC5_MAIN_CLK_GATE_FLD_PRBS_EN 0
`define DDRMC5_MAIN_CLK_GATE_FLD_PRBS_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CPLX_EN 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CPLX_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_ILECC_EN 2
`define DDRMC5_MAIN_CLK_GATE_FLD_ILECC_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN1_EN 3
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN1_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CAL_RD_DATA_EN 4
`define DDRMC5_MAIN_CLK_GATE_FLD_CAL_RD_DATA_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_DEBUG_EN 5
`define DDRMC5_MAIN_CLK_GATE_FLD_DEBUG_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CUST_PAT_EN 6
`define DDRMC5_MAIN_CLK_GATE_FLD_CUST_PAT_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_EDGE_DET_EN 7
`define DDRMC5_MAIN_CLK_GATE_FLD_EDGE_DET_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_ACC_EN 8
`define DDRMC5_MAIN_CLK_GATE_FLD_ACC_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CMPR_EN 9
`define DDRMC5_MAIN_CLK_GATE_FLD_CMPR_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_RESERVED 10
`define DDRMC5_MAIN_CLK_GATE_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU0_EN 11
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU0_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU1_EN 12
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU1_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU2_EN 13
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU2_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU3_EN 14
`define DDRMC5_MAIN_CLK_GATE_FLD_NSU3_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN0_DYN_GATE_DIS 15
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN0_DYN_GATE_DIS_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN1_DYN_GATE_DIS 16
`define DDRMC5_MAIN_CLK_GATE_FLD_CHAN1_DYN_GATE_DIS_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_NA_DYN_GATE_DIS 17
`define DDRMC5_MAIN_CLK_GATE_FLD_NA_DYN_GATE_DIS_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_DDRMC_EN 18
`define DDRMC5_MAIN_CLK_GATE_FLD_DDRMC_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_EN 19
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_XTS_EN 20
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_XTS_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_GCM_EN 21
`define DDRMC5_MAIN_CLK_GATE_FLD_CRYPTO_GCM_EN_WIDTH 1
`define DDRMC5_MAIN_CLK_GATE_FLD_RESERVED_1 31:22
`define DDRMC5_MAIN_CLK_GATE_FLD_RESERVED_1_WIDTH 10
`define DDRMC5_MAIN_CLK_GATE_WIDTH 22

/* ARBITER_CONFIG */
`define DDRMC5_MAIN_ARBITER_CONFIG_OFFSET 16'h91c
`define DDRMC5_MAIN_ARBITER_CONFIG_FLD_PRIORITY_SETTING 0
`define DDRMC5_MAIN_ARBITER_CONFIG_FLD_PRIORITY_SETTING_WIDTH 1
`define DDRMC5_MAIN_ARBITER_CONFIG_FLD_RESERVED 31:1
`define DDRMC5_MAIN_ARBITER_CONFIG_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_ARBITER_CONFIG_WIDTH 1

/* XPI_MRS_CONFIG */
`define DDRMC5_MAIN_XPI_MRS_CONFIG_OFFSET 16'h920
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_ENABLE 0
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_ENABLE_WIDTH 1
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_RESERVED 1
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_DDR5_BIT_SEL 2
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_DDR5_BIT_SEL_WIDTH 1
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_LP5_PHASE_SEL 5:3
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_LP5_PHASE_SEL_WIDTH 3
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_ERR_NIB_EN 15:6
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_ERR_NIB_EN_WIDTH 10
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_RESERVED_1 31:16
`define DDRMC5_MAIN_XPI_MRS_CONFIG_FLD_RESERVED_1_WIDTH 16
`define DDRMC5_MAIN_XPI_MRS_CONFIG_WIDTH 16

/* CPLX_PATTERN0 */
`define DDRMC5_MAIN_CPLX_PATTERN0_OFFSET 16'h924
`define DDRMC5_MAIN_CPLX_PATTERN0_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN0_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN0_WIDTH 16

/* CPLX_PATTERN1 */
`define DDRMC5_MAIN_CPLX_PATTERN1_OFFSET 16'h928
`define DDRMC5_MAIN_CPLX_PATTERN1_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN1_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN1_WIDTH 16

/* CPLX_PATTERN2 */
`define DDRMC5_MAIN_CPLX_PATTERN2_OFFSET 16'h92c
`define DDRMC5_MAIN_CPLX_PATTERN2_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN2_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN2_WIDTH 16

/* CPLX_PATTERN3 */
`define DDRMC5_MAIN_CPLX_PATTERN3_OFFSET 16'h930
`define DDRMC5_MAIN_CPLX_PATTERN3_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN3_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN3_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN3_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN3_WIDTH 16

/* CPLX_PATTERN4 */
`define DDRMC5_MAIN_CPLX_PATTERN4_OFFSET 16'h934
`define DDRMC5_MAIN_CPLX_PATTERN4_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN4_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN4_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN4_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN4_WIDTH 16

/* CPLX_PATTERN5 */
`define DDRMC5_MAIN_CPLX_PATTERN5_OFFSET 16'h938
`define DDRMC5_MAIN_CPLX_PATTERN5_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN5_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN5_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN5_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN5_WIDTH 16

/* CPLX_PATTERN6 */
`define DDRMC5_MAIN_CPLX_PATTERN6_OFFSET 16'h93c
`define DDRMC5_MAIN_CPLX_PATTERN6_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN6_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN6_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN6_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN6_WIDTH 16

/* CPLX_PATTERN7 */
`define DDRMC5_MAIN_CPLX_PATTERN7_OFFSET 16'h940
`define DDRMC5_MAIN_CPLX_PATTERN7_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN7_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN7_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN7_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN7_WIDTH 16

/* CPLX_PATTERN8 */
`define DDRMC5_MAIN_CPLX_PATTERN8_OFFSET 16'h944
`define DDRMC5_MAIN_CPLX_PATTERN8_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN8_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN8_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN8_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN8_WIDTH 16

/* CPLX_PATTERN9 */
`define DDRMC5_MAIN_CPLX_PATTERN9_OFFSET 16'h948
`define DDRMC5_MAIN_CPLX_PATTERN9_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN9_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN9_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN9_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN9_WIDTH 16

/* CPLX_PATTERN10 */
`define DDRMC5_MAIN_CPLX_PATTERN10_OFFSET 16'h94c
`define DDRMC5_MAIN_CPLX_PATTERN10_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN10_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN10_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN10_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN10_WIDTH 16

/* CPLX_PATTERN11 */
`define DDRMC5_MAIN_CPLX_PATTERN11_OFFSET 16'h950
`define DDRMC5_MAIN_CPLX_PATTERN11_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN11_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN11_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN11_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN11_WIDTH 16

/* CPLX_PATTERN12 */
`define DDRMC5_MAIN_CPLX_PATTERN12_OFFSET 16'h954
`define DDRMC5_MAIN_CPLX_PATTERN12_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN12_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN12_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN12_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN12_WIDTH 16

/* CPLX_PATTERN13 */
`define DDRMC5_MAIN_CPLX_PATTERN13_OFFSET 16'h958
`define DDRMC5_MAIN_CPLX_PATTERN13_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN13_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN13_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN13_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN13_WIDTH 16

/* CPLX_PATTERN14 */
`define DDRMC5_MAIN_CPLX_PATTERN14_OFFSET 16'h95c
`define DDRMC5_MAIN_CPLX_PATTERN14_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN14_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN14_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN14_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN14_WIDTH 16

/* CPLX_PATTERN15 */
`define DDRMC5_MAIN_CPLX_PATTERN15_OFFSET 16'h960
`define DDRMC5_MAIN_CPLX_PATTERN15_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN15_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN15_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN15_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN15_WIDTH 16

/* CPLX_PATTERN16 */
`define DDRMC5_MAIN_CPLX_PATTERN16_OFFSET 16'h964
`define DDRMC5_MAIN_CPLX_PATTERN16_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN16_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN16_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN16_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN16_WIDTH 16

/* CPLX_PATTERN17 */
`define DDRMC5_MAIN_CPLX_PATTERN17_OFFSET 16'h968
`define DDRMC5_MAIN_CPLX_PATTERN17_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN17_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN17_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN17_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN17_WIDTH 16

/* CPLX_PATTERN18 */
`define DDRMC5_MAIN_CPLX_PATTERN18_OFFSET 16'h96c
`define DDRMC5_MAIN_CPLX_PATTERN18_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN18_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN18_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN18_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN18_WIDTH 16

/* CPLX_PATTERN19 */
`define DDRMC5_MAIN_CPLX_PATTERN19_OFFSET 16'h970
`define DDRMC5_MAIN_CPLX_PATTERN19_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN19_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN19_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN19_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN19_WIDTH 16

/* CPLX_PATTERN20 */
`define DDRMC5_MAIN_CPLX_PATTERN20_OFFSET 16'h974
`define DDRMC5_MAIN_CPLX_PATTERN20_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN20_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN20_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN20_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN20_WIDTH 16

/* CPLX_PATTERN21 */
`define DDRMC5_MAIN_CPLX_PATTERN21_OFFSET 16'h978
`define DDRMC5_MAIN_CPLX_PATTERN21_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN21_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN21_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN21_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN21_WIDTH 16

/* CPLX_PATTERN22 */
`define DDRMC5_MAIN_CPLX_PATTERN22_OFFSET 16'h97c
`define DDRMC5_MAIN_CPLX_PATTERN22_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN22_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN22_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN22_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN22_WIDTH 16

/* CPLX_PATTERN23 */
`define DDRMC5_MAIN_CPLX_PATTERN23_OFFSET 16'h980
`define DDRMC5_MAIN_CPLX_PATTERN23_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN23_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN23_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN23_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN23_WIDTH 16

/* CPLX_PATTERN24 */
`define DDRMC5_MAIN_CPLX_PATTERN24_OFFSET 16'h984
`define DDRMC5_MAIN_CPLX_PATTERN24_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN24_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN24_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN24_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN24_WIDTH 16

/* CPLX_PATTERN25 */
`define DDRMC5_MAIN_CPLX_PATTERN25_OFFSET 16'h988
`define DDRMC5_MAIN_CPLX_PATTERN25_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN25_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN25_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN25_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN25_WIDTH 16

/* CPLX_PATTERN26 */
`define DDRMC5_MAIN_CPLX_PATTERN26_OFFSET 16'h98c
`define DDRMC5_MAIN_CPLX_PATTERN26_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN26_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN26_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN26_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN26_WIDTH 16

/* CPLX_PATTERN27 */
`define DDRMC5_MAIN_CPLX_PATTERN27_OFFSET 16'h990
`define DDRMC5_MAIN_CPLX_PATTERN27_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN27_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN27_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN27_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN27_WIDTH 16

/* CPLX_PATTERN28 */
`define DDRMC5_MAIN_CPLX_PATTERN28_OFFSET 16'h994
`define DDRMC5_MAIN_CPLX_PATTERN28_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN28_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN28_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN28_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN28_WIDTH 16

/* CPLX_PATTERN29 */
`define DDRMC5_MAIN_CPLX_PATTERN29_OFFSET 16'h998
`define DDRMC5_MAIN_CPLX_PATTERN29_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN29_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN29_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN29_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN29_WIDTH 16

/* CPLX_PATTERN30 */
`define DDRMC5_MAIN_CPLX_PATTERN30_OFFSET 16'h99c
`define DDRMC5_MAIN_CPLX_PATTERN30_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN30_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN30_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN30_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN30_WIDTH 16

/* CPLX_PATTERN31 */
`define DDRMC5_MAIN_CPLX_PATTERN31_OFFSET 16'h9a0
`define DDRMC5_MAIN_CPLX_PATTERN31_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN31_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN31_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN31_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN31_WIDTH 16

/* CPLX_PATTERN32 */
`define DDRMC5_MAIN_CPLX_PATTERN32_OFFSET 16'h9a4
`define DDRMC5_MAIN_CPLX_PATTERN32_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN32_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN32_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN32_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN32_WIDTH 16

/* CPLX_PATTERN33 */
`define DDRMC5_MAIN_CPLX_PATTERN33_OFFSET 16'h9a8
`define DDRMC5_MAIN_CPLX_PATTERN33_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN33_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN33_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN33_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN33_WIDTH 16

/* CPLX_PATTERN34 */
`define DDRMC5_MAIN_CPLX_PATTERN34_OFFSET 16'h9ac
`define DDRMC5_MAIN_CPLX_PATTERN34_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN34_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN34_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN34_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN34_WIDTH 16

/* CPLX_PATTERN35 */
`define DDRMC5_MAIN_CPLX_PATTERN35_OFFSET 16'h9b0
`define DDRMC5_MAIN_CPLX_PATTERN35_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN35_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN35_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN35_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN35_WIDTH 16

/* CPLX_PATTERN36 */
`define DDRMC5_MAIN_CPLX_PATTERN36_OFFSET 16'h9b4
`define DDRMC5_MAIN_CPLX_PATTERN36_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN36_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN36_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN36_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN36_WIDTH 16

/* CPLX_PATTERN37 */
`define DDRMC5_MAIN_CPLX_PATTERN37_OFFSET 16'h9b8
`define DDRMC5_MAIN_CPLX_PATTERN37_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN37_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN37_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN37_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN37_WIDTH 16

/* CPLX_PATTERN38 */
`define DDRMC5_MAIN_CPLX_PATTERN38_OFFSET 16'h9bc
`define DDRMC5_MAIN_CPLX_PATTERN38_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN38_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN38_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN38_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN38_WIDTH 16

/* CPLX_PATTERN39 */
`define DDRMC5_MAIN_CPLX_PATTERN39_OFFSET 16'h9c0
`define DDRMC5_MAIN_CPLX_PATTERN39_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN39_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN39_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN39_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN39_WIDTH 16

/* CPLX_PATTERN40 */
`define DDRMC5_MAIN_CPLX_PATTERN40_OFFSET 16'h9c4
`define DDRMC5_MAIN_CPLX_PATTERN40_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN40_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN40_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN40_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN40_WIDTH 16

/* CPLX_PATTERN41 */
`define DDRMC5_MAIN_CPLX_PATTERN41_OFFSET 16'h9c8
`define DDRMC5_MAIN_CPLX_PATTERN41_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN41_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN41_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN41_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN41_WIDTH 16

/* CPLX_PATTERN42 */
`define DDRMC5_MAIN_CPLX_PATTERN42_OFFSET 16'h9cc
`define DDRMC5_MAIN_CPLX_PATTERN42_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN42_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN42_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN42_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN42_WIDTH 16

/* CPLX_PATTERN43 */
`define DDRMC5_MAIN_CPLX_PATTERN43_OFFSET 16'h9d0
`define DDRMC5_MAIN_CPLX_PATTERN43_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN43_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN43_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN43_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN43_WIDTH 16

/* CPLX_PATTERN44 */
`define DDRMC5_MAIN_CPLX_PATTERN44_OFFSET 16'h9d4
`define DDRMC5_MAIN_CPLX_PATTERN44_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN44_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN44_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN44_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN44_WIDTH 16

/* CPLX_PATTERN45 */
`define DDRMC5_MAIN_CPLX_PATTERN45_OFFSET 16'h9d8
`define DDRMC5_MAIN_CPLX_PATTERN45_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN45_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN45_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN45_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN45_WIDTH 16

/* CPLX_PATTERN46 */
`define DDRMC5_MAIN_CPLX_PATTERN46_OFFSET 16'h9dc
`define DDRMC5_MAIN_CPLX_PATTERN46_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN46_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN46_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN46_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN46_WIDTH 16

/* CPLX_PATTERN47 */
`define DDRMC5_MAIN_CPLX_PATTERN47_OFFSET 16'h9e0
`define DDRMC5_MAIN_CPLX_PATTERN47_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN47_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN47_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN47_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN47_WIDTH 16

/* CPLX_PATTERN48 */
`define DDRMC5_MAIN_CPLX_PATTERN48_OFFSET 16'h9e4
`define DDRMC5_MAIN_CPLX_PATTERN48_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN48_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN48_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN48_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN48_WIDTH 16

/* CPLX_PATTERN49 */
`define DDRMC5_MAIN_CPLX_PATTERN49_OFFSET 16'h9e8
`define DDRMC5_MAIN_CPLX_PATTERN49_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN49_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN49_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN49_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN49_WIDTH 16

/* CPLX_PATTERN50 */
`define DDRMC5_MAIN_CPLX_PATTERN50_OFFSET 16'h9ec
`define DDRMC5_MAIN_CPLX_PATTERN50_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN50_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN50_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN50_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN50_WIDTH 16

/* CPLX_PATTERN51 */
`define DDRMC5_MAIN_CPLX_PATTERN51_OFFSET 16'h9f0
`define DDRMC5_MAIN_CPLX_PATTERN51_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN51_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN51_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN51_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN51_WIDTH 16

/* CPLX_PATTERN52 */
`define DDRMC5_MAIN_CPLX_PATTERN52_OFFSET 16'h9f4
`define DDRMC5_MAIN_CPLX_PATTERN52_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN52_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN52_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN52_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN52_WIDTH 16

/* CPLX_PATTERN53 */
`define DDRMC5_MAIN_CPLX_PATTERN53_OFFSET 16'h9f8
`define DDRMC5_MAIN_CPLX_PATTERN53_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN53_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN53_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN53_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN53_WIDTH 16

/* CPLX_PATTERN54 */
`define DDRMC5_MAIN_CPLX_PATTERN54_OFFSET 16'h9fc
`define DDRMC5_MAIN_CPLX_PATTERN54_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN54_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN54_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN54_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN54_WIDTH 16

/* CPLX_PATTERN55 */
`define DDRMC5_MAIN_CPLX_PATTERN55_OFFSET 16'ha00
`define DDRMC5_MAIN_CPLX_PATTERN55_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN55_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN55_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN55_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN55_WIDTH 16

/* CPLX_PATTERN56 */
`define DDRMC5_MAIN_CPLX_PATTERN56_OFFSET 16'ha04
`define DDRMC5_MAIN_CPLX_PATTERN56_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN56_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN56_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN56_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN56_WIDTH 16

/* CPLX_PATTERN57 */
`define DDRMC5_MAIN_CPLX_PATTERN57_OFFSET 16'ha08
`define DDRMC5_MAIN_CPLX_PATTERN57_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN57_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN57_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN57_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN57_WIDTH 16

/* CPLX_PATTERN58 */
`define DDRMC5_MAIN_CPLX_PATTERN58_OFFSET 16'ha0c
`define DDRMC5_MAIN_CPLX_PATTERN58_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN58_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN58_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN58_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN58_WIDTH 16

/* CPLX_PATTERN59 */
`define DDRMC5_MAIN_CPLX_PATTERN59_OFFSET 16'ha10
`define DDRMC5_MAIN_CPLX_PATTERN59_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN59_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN59_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN59_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN59_WIDTH 16

/* CPLX_PATTERN60 */
`define DDRMC5_MAIN_CPLX_PATTERN60_OFFSET 16'ha14
`define DDRMC5_MAIN_CPLX_PATTERN60_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN60_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN60_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN60_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN60_WIDTH 16

/* CPLX_PATTERN61 */
`define DDRMC5_MAIN_CPLX_PATTERN61_OFFSET 16'ha18
`define DDRMC5_MAIN_CPLX_PATTERN61_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN61_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN61_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN61_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN61_WIDTH 16

/* CPLX_PATTERN62 */
`define DDRMC5_MAIN_CPLX_PATTERN62_OFFSET 16'ha1c
`define DDRMC5_MAIN_CPLX_PATTERN62_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN62_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN62_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN62_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN62_WIDTH 16

/* CPLX_PATTERN63 */
`define DDRMC5_MAIN_CPLX_PATTERN63_OFFSET 16'ha20
`define DDRMC5_MAIN_CPLX_PATTERN63_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN63_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN63_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN63_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN63_WIDTH 16

/* CPLX_PATTERN64 */
`define DDRMC5_MAIN_CPLX_PATTERN64_OFFSET 16'ha24
`define DDRMC5_MAIN_CPLX_PATTERN64_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN64_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN64_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN64_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN64_WIDTH 16

/* CPLX_PATTERN65 */
`define DDRMC5_MAIN_CPLX_PATTERN65_OFFSET 16'ha28
`define DDRMC5_MAIN_CPLX_PATTERN65_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN65_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN65_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN65_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN65_WIDTH 16

/* CPLX_PATTERN66 */
`define DDRMC5_MAIN_CPLX_PATTERN66_OFFSET 16'ha2c
`define DDRMC5_MAIN_CPLX_PATTERN66_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN66_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN66_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN66_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN66_WIDTH 16

/* CPLX_PATTERN67 */
`define DDRMC5_MAIN_CPLX_PATTERN67_OFFSET 16'ha30
`define DDRMC5_MAIN_CPLX_PATTERN67_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN67_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN67_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN67_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN67_WIDTH 16

/* CPLX_PATTERN68 */
`define DDRMC5_MAIN_CPLX_PATTERN68_OFFSET 16'ha34
`define DDRMC5_MAIN_CPLX_PATTERN68_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN68_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN68_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN68_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN68_WIDTH 16

/* CPLX_PATTERN69 */
`define DDRMC5_MAIN_CPLX_PATTERN69_OFFSET 16'ha38
`define DDRMC5_MAIN_CPLX_PATTERN69_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN69_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN69_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN69_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN69_WIDTH 16

/* CPLX_PATTERN70 */
`define DDRMC5_MAIN_CPLX_PATTERN70_OFFSET 16'ha3c
`define DDRMC5_MAIN_CPLX_PATTERN70_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN70_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN70_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN70_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN70_WIDTH 16

/* CPLX_PATTERN71 */
`define DDRMC5_MAIN_CPLX_PATTERN71_OFFSET 16'ha40
`define DDRMC5_MAIN_CPLX_PATTERN71_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN71_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN71_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN71_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN71_WIDTH 16

/* CPLX_PATTERN72 */
`define DDRMC5_MAIN_CPLX_PATTERN72_OFFSET 16'ha44
`define DDRMC5_MAIN_CPLX_PATTERN72_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN72_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN72_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN72_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN72_WIDTH 16

/* CPLX_PATTERN73 */
`define DDRMC5_MAIN_CPLX_PATTERN73_OFFSET 16'ha48
`define DDRMC5_MAIN_CPLX_PATTERN73_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN73_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN73_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN73_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN73_WIDTH 16

/* CPLX_PATTERN74 */
`define DDRMC5_MAIN_CPLX_PATTERN74_OFFSET 16'ha4c
`define DDRMC5_MAIN_CPLX_PATTERN74_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN74_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN74_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN74_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN74_WIDTH 16

/* CPLX_PATTERN75 */
`define DDRMC5_MAIN_CPLX_PATTERN75_OFFSET 16'ha50
`define DDRMC5_MAIN_CPLX_PATTERN75_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN75_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN75_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN75_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN75_WIDTH 16

/* CPLX_PATTERN76 */
`define DDRMC5_MAIN_CPLX_PATTERN76_OFFSET 16'ha54
`define DDRMC5_MAIN_CPLX_PATTERN76_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN76_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN76_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN76_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN76_WIDTH 16

/* CPLX_PATTERN77 */
`define DDRMC5_MAIN_CPLX_PATTERN77_OFFSET 16'ha58
`define DDRMC5_MAIN_CPLX_PATTERN77_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN77_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN77_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN77_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN77_WIDTH 16

/* CPLX_PATTERN78 */
`define DDRMC5_MAIN_CPLX_PATTERN78_OFFSET 16'ha5c
`define DDRMC5_MAIN_CPLX_PATTERN78_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN78_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN78_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN78_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN78_WIDTH 16

/* CPLX_PATTERN79 */
`define DDRMC5_MAIN_CPLX_PATTERN79_OFFSET 16'ha60
`define DDRMC5_MAIN_CPLX_PATTERN79_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN79_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN79_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN79_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN79_WIDTH 16

/* CPLX_PATTERN80 */
`define DDRMC5_MAIN_CPLX_PATTERN80_OFFSET 16'ha64
`define DDRMC5_MAIN_CPLX_PATTERN80_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN80_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN80_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN80_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN80_WIDTH 16

/* CPLX_PATTERN81 */
`define DDRMC5_MAIN_CPLX_PATTERN81_OFFSET 16'ha68
`define DDRMC5_MAIN_CPLX_PATTERN81_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN81_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN81_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN81_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN81_WIDTH 16

/* CPLX_PATTERN82 */
`define DDRMC5_MAIN_CPLX_PATTERN82_OFFSET 16'ha6c
`define DDRMC5_MAIN_CPLX_PATTERN82_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN82_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN82_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN82_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN82_WIDTH 16

/* CPLX_PATTERN83 */
`define DDRMC5_MAIN_CPLX_PATTERN83_OFFSET 16'ha70
`define DDRMC5_MAIN_CPLX_PATTERN83_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN83_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN83_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN83_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN83_WIDTH 16

/* CPLX_PATTERN84 */
`define DDRMC5_MAIN_CPLX_PATTERN84_OFFSET 16'ha74
`define DDRMC5_MAIN_CPLX_PATTERN84_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN84_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN84_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN84_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN84_WIDTH 16

/* CPLX_PATTERN85 */
`define DDRMC5_MAIN_CPLX_PATTERN85_OFFSET 16'ha78
`define DDRMC5_MAIN_CPLX_PATTERN85_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN85_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN85_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN85_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN85_WIDTH 16

/* CPLX_PATTERN86 */
`define DDRMC5_MAIN_CPLX_PATTERN86_OFFSET 16'ha7c
`define DDRMC5_MAIN_CPLX_PATTERN86_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN86_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN86_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN86_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN86_WIDTH 16

/* CPLX_PATTERN87 */
`define DDRMC5_MAIN_CPLX_PATTERN87_OFFSET 16'ha80
`define DDRMC5_MAIN_CPLX_PATTERN87_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN87_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN87_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN87_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN87_WIDTH 16

/* CPLX_PATTERN88 */
`define DDRMC5_MAIN_CPLX_PATTERN88_OFFSET 16'ha84
`define DDRMC5_MAIN_CPLX_PATTERN88_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN88_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN88_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN88_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN88_WIDTH 16

/* CPLX_PATTERN89 */
`define DDRMC5_MAIN_CPLX_PATTERN89_OFFSET 16'ha88
`define DDRMC5_MAIN_CPLX_PATTERN89_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN89_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN89_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN89_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN89_WIDTH 16

/* CPLX_PATTERN90 */
`define DDRMC5_MAIN_CPLX_PATTERN90_OFFSET 16'ha8c
`define DDRMC5_MAIN_CPLX_PATTERN90_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN90_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN90_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN90_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN90_WIDTH 16

/* CPLX_PATTERN91 */
`define DDRMC5_MAIN_CPLX_PATTERN91_OFFSET 16'ha90
`define DDRMC5_MAIN_CPLX_PATTERN91_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN91_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN91_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN91_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN91_WIDTH 16

/* CPLX_PATTERN92 */
`define DDRMC5_MAIN_CPLX_PATTERN92_OFFSET 16'ha94
`define DDRMC5_MAIN_CPLX_PATTERN92_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN92_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN92_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN92_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN92_WIDTH 16

/* CPLX_PATTERN93 */
`define DDRMC5_MAIN_CPLX_PATTERN93_OFFSET 16'ha98
`define DDRMC5_MAIN_CPLX_PATTERN93_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN93_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN93_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN93_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN93_WIDTH 16

/* CPLX_PATTERN94 */
`define DDRMC5_MAIN_CPLX_PATTERN94_OFFSET 16'ha9c
`define DDRMC5_MAIN_CPLX_PATTERN94_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN94_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN94_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN94_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN94_WIDTH 16

/* CPLX_PATTERN95 */
`define DDRMC5_MAIN_CPLX_PATTERN95_OFFSET 16'haa0
`define DDRMC5_MAIN_CPLX_PATTERN95_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN95_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN95_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN95_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN95_WIDTH 16

/* CPLX_PATTERN96 */
`define DDRMC5_MAIN_CPLX_PATTERN96_OFFSET 16'haa4
`define DDRMC5_MAIN_CPLX_PATTERN96_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN96_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN96_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN96_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN96_WIDTH 16

/* CPLX_PATTERN97 */
`define DDRMC5_MAIN_CPLX_PATTERN97_OFFSET 16'haa8
`define DDRMC5_MAIN_CPLX_PATTERN97_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN97_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN97_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN97_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN97_WIDTH 16

/* CPLX_PATTERN98 */
`define DDRMC5_MAIN_CPLX_PATTERN98_OFFSET 16'haac
`define DDRMC5_MAIN_CPLX_PATTERN98_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN98_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN98_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN98_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN98_WIDTH 16

/* CPLX_PATTERN99 */
`define DDRMC5_MAIN_CPLX_PATTERN99_OFFSET 16'hab0
`define DDRMC5_MAIN_CPLX_PATTERN99_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN99_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN99_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN99_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN99_WIDTH 16

/* CPLX_PATTERN100 */
`define DDRMC5_MAIN_CPLX_PATTERN100_OFFSET 16'hab4
`define DDRMC5_MAIN_CPLX_PATTERN100_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN100_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN100_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN100_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN100_WIDTH 16

/* CPLX_PATTERN101 */
`define DDRMC5_MAIN_CPLX_PATTERN101_OFFSET 16'hab8
`define DDRMC5_MAIN_CPLX_PATTERN101_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN101_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN101_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN101_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN101_WIDTH 16

/* CPLX_PATTERN102 */
`define DDRMC5_MAIN_CPLX_PATTERN102_OFFSET 16'habc
`define DDRMC5_MAIN_CPLX_PATTERN102_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN102_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN102_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN102_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN102_WIDTH 16

/* CPLX_PATTERN103 */
`define DDRMC5_MAIN_CPLX_PATTERN103_OFFSET 16'hac0
`define DDRMC5_MAIN_CPLX_PATTERN103_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN103_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN103_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN103_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN103_WIDTH 16

/* CPLX_PATTERN104 */
`define DDRMC5_MAIN_CPLX_PATTERN104_OFFSET 16'hac4
`define DDRMC5_MAIN_CPLX_PATTERN104_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN104_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN104_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN104_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN104_WIDTH 16

/* CPLX_PATTERN105 */
`define DDRMC5_MAIN_CPLX_PATTERN105_OFFSET 16'hac8
`define DDRMC5_MAIN_CPLX_PATTERN105_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN105_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN105_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN105_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN105_WIDTH 16

/* CPLX_PATTERN106 */
`define DDRMC5_MAIN_CPLX_PATTERN106_OFFSET 16'hacc
`define DDRMC5_MAIN_CPLX_PATTERN106_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN106_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN106_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN106_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN106_WIDTH 16

/* CPLX_PATTERN107 */
`define DDRMC5_MAIN_CPLX_PATTERN107_OFFSET 16'had0
`define DDRMC5_MAIN_CPLX_PATTERN107_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN107_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN107_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN107_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN107_WIDTH 16

/* CPLX_PATTERN108 */
`define DDRMC5_MAIN_CPLX_PATTERN108_OFFSET 16'had4
`define DDRMC5_MAIN_CPLX_PATTERN108_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN108_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN108_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN108_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN108_WIDTH 16

/* CPLX_PATTERN109 */
`define DDRMC5_MAIN_CPLX_PATTERN109_OFFSET 16'had8
`define DDRMC5_MAIN_CPLX_PATTERN109_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN109_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN109_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN109_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN109_WIDTH 16

/* CPLX_PATTERN110 */
`define DDRMC5_MAIN_CPLX_PATTERN110_OFFSET 16'hadc
`define DDRMC5_MAIN_CPLX_PATTERN110_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN110_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN110_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN110_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN110_WIDTH 16

/* CPLX_PATTERN111 */
`define DDRMC5_MAIN_CPLX_PATTERN111_OFFSET 16'hae0
`define DDRMC5_MAIN_CPLX_PATTERN111_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN111_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN111_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN111_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN111_WIDTH 16

/* CPLX_PATTERN112 */
`define DDRMC5_MAIN_CPLX_PATTERN112_OFFSET 16'hae4
`define DDRMC5_MAIN_CPLX_PATTERN112_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN112_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN112_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN112_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN112_WIDTH 16

/* CPLX_PATTERN113 */
`define DDRMC5_MAIN_CPLX_PATTERN113_OFFSET 16'hae8
`define DDRMC5_MAIN_CPLX_PATTERN113_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN113_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN113_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN113_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN113_WIDTH 16

/* CPLX_PATTERN114 */
`define DDRMC5_MAIN_CPLX_PATTERN114_OFFSET 16'haec
`define DDRMC5_MAIN_CPLX_PATTERN114_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN114_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN114_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN114_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN114_WIDTH 16

/* CPLX_PATTERN115 */
`define DDRMC5_MAIN_CPLX_PATTERN115_OFFSET 16'haf0
`define DDRMC5_MAIN_CPLX_PATTERN115_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN115_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN115_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN115_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN115_WIDTH 16

/* CPLX_PATTERN116 */
`define DDRMC5_MAIN_CPLX_PATTERN116_OFFSET 16'haf4
`define DDRMC5_MAIN_CPLX_PATTERN116_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN116_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN116_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN116_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN116_WIDTH 16

/* CPLX_PATTERN117 */
`define DDRMC5_MAIN_CPLX_PATTERN117_OFFSET 16'haf8
`define DDRMC5_MAIN_CPLX_PATTERN117_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN117_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN117_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN117_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN117_WIDTH 16

/* CPLX_PATTERN118 */
`define DDRMC5_MAIN_CPLX_PATTERN118_OFFSET 16'hafc
`define DDRMC5_MAIN_CPLX_PATTERN118_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN118_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN118_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN118_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN118_WIDTH 16

/* CPLX_PATTERN119 */
`define DDRMC5_MAIN_CPLX_PATTERN119_OFFSET 16'hb00
`define DDRMC5_MAIN_CPLX_PATTERN119_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN119_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN119_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN119_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN119_WIDTH 16

/* CPLX_PATTERN120 */
`define DDRMC5_MAIN_CPLX_PATTERN120_OFFSET 16'hb04
`define DDRMC5_MAIN_CPLX_PATTERN120_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN120_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN120_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN120_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN120_WIDTH 16

/* CPLX_PATTERN121 */
`define DDRMC5_MAIN_CPLX_PATTERN121_OFFSET 16'hb08
`define DDRMC5_MAIN_CPLX_PATTERN121_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN121_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN121_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN121_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN121_WIDTH 16

/* CPLX_PATTERN122 */
`define DDRMC5_MAIN_CPLX_PATTERN122_OFFSET 16'hb0c
`define DDRMC5_MAIN_CPLX_PATTERN122_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN122_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN122_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN122_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN122_WIDTH 16

/* CPLX_PATTERN123 */
`define DDRMC5_MAIN_CPLX_PATTERN123_OFFSET 16'hb10
`define DDRMC5_MAIN_CPLX_PATTERN123_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN123_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN123_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN123_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN123_WIDTH 16

/* CPLX_PATTERN124 */
`define DDRMC5_MAIN_CPLX_PATTERN124_OFFSET 16'hb14
`define DDRMC5_MAIN_CPLX_PATTERN124_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN124_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN124_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN124_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN124_WIDTH 16

/* CPLX_PATTERN125 */
`define DDRMC5_MAIN_CPLX_PATTERN125_OFFSET 16'hb18
`define DDRMC5_MAIN_CPLX_PATTERN125_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN125_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN125_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN125_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN125_WIDTH 16

/* CPLX_PATTERN126 */
`define DDRMC5_MAIN_CPLX_PATTERN126_OFFSET 16'hb1c
`define DDRMC5_MAIN_CPLX_PATTERN126_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN126_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN126_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN126_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN126_WIDTH 16

/* CPLX_PATTERN127 */
`define DDRMC5_MAIN_CPLX_PATTERN127_OFFSET 16'hb20
`define DDRMC5_MAIN_CPLX_PATTERN127_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN127_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN127_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN127_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN127_WIDTH 16

/* CPLX_PATTERN128 */
`define DDRMC5_MAIN_CPLX_PATTERN128_OFFSET 16'hb24
`define DDRMC5_MAIN_CPLX_PATTERN128_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN128_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN128_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN128_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN128_WIDTH 16

/* CPLX_PATTERN129 */
`define DDRMC5_MAIN_CPLX_PATTERN129_OFFSET 16'hb28
`define DDRMC5_MAIN_CPLX_PATTERN129_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN129_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN129_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN129_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN129_WIDTH 16

/* CPLX_PATTERN130 */
`define DDRMC5_MAIN_CPLX_PATTERN130_OFFSET 16'hb2c
`define DDRMC5_MAIN_CPLX_PATTERN130_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN130_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN130_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN130_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN130_WIDTH 16

/* CPLX_PATTERN131 */
`define DDRMC5_MAIN_CPLX_PATTERN131_OFFSET 16'hb30
`define DDRMC5_MAIN_CPLX_PATTERN131_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN131_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN131_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN131_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN131_WIDTH 16

/* CPLX_PATTERN132 */
`define DDRMC5_MAIN_CPLX_PATTERN132_OFFSET 16'hb34
`define DDRMC5_MAIN_CPLX_PATTERN132_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN132_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN132_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN132_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN132_WIDTH 16

/* CPLX_PATTERN133 */
`define DDRMC5_MAIN_CPLX_PATTERN133_OFFSET 16'hb38
`define DDRMC5_MAIN_CPLX_PATTERN133_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN133_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN133_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN133_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN133_WIDTH 16

/* CPLX_PATTERN134 */
`define DDRMC5_MAIN_CPLX_PATTERN134_OFFSET 16'hb3c
`define DDRMC5_MAIN_CPLX_PATTERN134_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN134_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN134_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN134_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN134_WIDTH 16

/* CPLX_PATTERN135 */
`define DDRMC5_MAIN_CPLX_PATTERN135_OFFSET 16'hb40
`define DDRMC5_MAIN_CPLX_PATTERN135_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN135_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN135_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN135_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN135_WIDTH 16

/* CPLX_PATTERN136 */
`define DDRMC5_MAIN_CPLX_PATTERN136_OFFSET 16'hb44
`define DDRMC5_MAIN_CPLX_PATTERN136_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN136_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN136_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN136_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN136_WIDTH 16

/* CPLX_PATTERN137 */
`define DDRMC5_MAIN_CPLX_PATTERN137_OFFSET 16'hb48
`define DDRMC5_MAIN_CPLX_PATTERN137_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN137_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN137_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN137_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN137_WIDTH 16

/* CPLX_PATTERN138 */
`define DDRMC5_MAIN_CPLX_PATTERN138_OFFSET 16'hb4c
`define DDRMC5_MAIN_CPLX_PATTERN138_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN138_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN138_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN138_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN138_WIDTH 16

/* CPLX_PATTERN139 */
`define DDRMC5_MAIN_CPLX_PATTERN139_OFFSET 16'hb50
`define DDRMC5_MAIN_CPLX_PATTERN139_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN139_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN139_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN139_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN139_WIDTH 16

/* CPLX_PATTERN140 */
`define DDRMC5_MAIN_CPLX_PATTERN140_OFFSET 16'hb54
`define DDRMC5_MAIN_CPLX_PATTERN140_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN140_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN140_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN140_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN140_WIDTH 16

/* CPLX_PATTERN141 */
`define DDRMC5_MAIN_CPLX_PATTERN141_OFFSET 16'hb58
`define DDRMC5_MAIN_CPLX_PATTERN141_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN141_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN141_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN141_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN141_WIDTH 16

/* CPLX_PATTERN142 */
`define DDRMC5_MAIN_CPLX_PATTERN142_OFFSET 16'hb5c
`define DDRMC5_MAIN_CPLX_PATTERN142_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN142_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN142_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN142_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN142_WIDTH 16

/* CPLX_PATTERN143 */
`define DDRMC5_MAIN_CPLX_PATTERN143_OFFSET 16'hb60
`define DDRMC5_MAIN_CPLX_PATTERN143_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN143_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN143_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN143_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN143_WIDTH 16

/* CPLX_PATTERN144 */
`define DDRMC5_MAIN_CPLX_PATTERN144_OFFSET 16'hb64
`define DDRMC5_MAIN_CPLX_PATTERN144_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN144_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN144_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN144_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN144_WIDTH 16

/* CPLX_PATTERN145 */
`define DDRMC5_MAIN_CPLX_PATTERN145_OFFSET 16'hb68
`define DDRMC5_MAIN_CPLX_PATTERN145_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN145_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN145_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN145_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN145_WIDTH 16

/* CPLX_PATTERN146 */
`define DDRMC5_MAIN_CPLX_PATTERN146_OFFSET 16'hb6c
`define DDRMC5_MAIN_CPLX_PATTERN146_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN146_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN146_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN146_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN146_WIDTH 16

/* CPLX_PATTERN147 */
`define DDRMC5_MAIN_CPLX_PATTERN147_OFFSET 16'hb70
`define DDRMC5_MAIN_CPLX_PATTERN147_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN147_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN147_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN147_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN147_WIDTH 16

/* CPLX_PATTERN148 */
`define DDRMC5_MAIN_CPLX_PATTERN148_OFFSET 16'hb74
`define DDRMC5_MAIN_CPLX_PATTERN148_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN148_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN148_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN148_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN148_WIDTH 16

/* CPLX_PATTERN149 */
`define DDRMC5_MAIN_CPLX_PATTERN149_OFFSET 16'hb78
`define DDRMC5_MAIN_CPLX_PATTERN149_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN149_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN149_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN149_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN149_WIDTH 16

/* CPLX_PATTERN150 */
`define DDRMC5_MAIN_CPLX_PATTERN150_OFFSET 16'hb7c
`define DDRMC5_MAIN_CPLX_PATTERN150_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN150_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN150_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN150_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN150_WIDTH 16

/* CPLX_PATTERN151 */
`define DDRMC5_MAIN_CPLX_PATTERN151_OFFSET 16'hb80
`define DDRMC5_MAIN_CPLX_PATTERN151_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN151_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN151_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN151_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN151_WIDTH 16

/* CPLX_PATTERN152 */
`define DDRMC5_MAIN_CPLX_PATTERN152_OFFSET 16'hb84
`define DDRMC5_MAIN_CPLX_PATTERN152_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN152_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN152_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN152_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN152_WIDTH 16

/* CPLX_PATTERN153 */
`define DDRMC5_MAIN_CPLX_PATTERN153_OFFSET 16'hb88
`define DDRMC5_MAIN_CPLX_PATTERN153_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN153_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN153_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN153_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN153_WIDTH 16

/* CPLX_PATTERN154 */
`define DDRMC5_MAIN_CPLX_PATTERN154_OFFSET 16'hb8c
`define DDRMC5_MAIN_CPLX_PATTERN154_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN154_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN154_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN154_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN154_WIDTH 16

/* CPLX_PATTERN155 */
`define DDRMC5_MAIN_CPLX_PATTERN155_OFFSET 16'hb90
`define DDRMC5_MAIN_CPLX_PATTERN155_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN155_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN155_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN155_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN155_WIDTH 16

/* CPLX_PATTERN156 */
`define DDRMC5_MAIN_CPLX_PATTERN156_OFFSET 16'hb94
`define DDRMC5_MAIN_CPLX_PATTERN156_FLD_VAL 15:0
`define DDRMC5_MAIN_CPLX_PATTERN156_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN156_FLD_RESERVED 31:16
`define DDRMC5_MAIN_CPLX_PATTERN156_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_CPLX_PATTERN156_WIDTH 16

/* CPLX_CONFIG2 */
`define DDRMC5_MAIN_CPLX_CONFIG2_OFFSET 16'hb98
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_WR_GAP_TIMER_VAL 4:0
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_WR_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RD_GAP_TIMER_VAL 9:5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RD_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_WR_BURST_GAP_TIMER_VAL 14:10
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_WR_BURST_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RD_BURST_GAP_TIMER_VAL 19:15
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RD_BURST_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_TWOBGBITSMODE_GAP_TIMER_VAL 24:20
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_TWOBGBITSMODE_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RESERVED 31:25
`define DDRMC5_MAIN_CPLX_CONFIG2_FLD_RESERVED_WIDTH 7
`define DDRMC5_MAIN_CPLX_CONFIG2_WIDTH 25

/* CPLX_BURST_ARRAY0 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_OFFSET 16'hb9c
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY0_WIDTH 5

/* CPLX_BURST_ARRAY1 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_OFFSET 16'hba0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY1_WIDTH 5

/* CPLX_BURST_ARRAY2 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_OFFSET 16'hba4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY2_WIDTH 5

/* CPLX_BURST_ARRAY3 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_OFFSET 16'hba8
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY3_WIDTH 5

/* CPLX_BURST_ARRAY4 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_OFFSET 16'hbac
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY4_WIDTH 5

/* CPLX_BURST_ARRAY5 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_OFFSET 16'hbb0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY5_WIDTH 5

/* CPLX_BURST_ARRAY6 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_OFFSET 16'hbb4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY6_WIDTH 5

/* CPLX_BURST_ARRAY7 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_OFFSET 16'hbb8
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY7_WIDTH 5

/* CPLX_BURST_ARRAY8 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_OFFSET 16'hbbc
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY8_WIDTH 5

/* CPLX_BURST_ARRAY9 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_OFFSET 16'hbc0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY9_WIDTH 5

/* CPLX_BURST_ARRAY10 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_OFFSET 16'hbc4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY10_WIDTH 5

/* CPLX_BURST_ARRAY11 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_OFFSET 16'hbc8
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY11_WIDTH 5

/* CPLX_BURST_ARRAY12 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_OFFSET 16'hbcc
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY12_WIDTH 5

/* CPLX_BURST_ARRAY13 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_OFFSET 16'hbd0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY13_WIDTH 5

/* CPLX_BURST_ARRAY14 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_OFFSET 16'hbd4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY14_WIDTH 5

/* CPLX_BURST_ARRAY15 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_OFFSET 16'hbd8
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY15_WIDTH 5

/* CPLX_BURST_ARRAY16 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_OFFSET 16'hbdc
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY16_WIDTH 5

/* CPLX_BURST_ARRAY17 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_OFFSET 16'hbe0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY17_WIDTH 5

/* CPLX_BURST_ARRAY18 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_OFFSET 16'hbe4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY18_WIDTH 5

/* CPLX_BURST_ARRAY19 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_OFFSET 16'hbe8
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY19_WIDTH 5

/* CPLX_BURST_ARRAY20 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_OFFSET 16'hbec
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY20_WIDTH 5

/* CPLX_BURST_ARRAY21 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_OFFSET 16'hbf0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY21_WIDTH 5

/* CPLX_BURST_ARRAY22 */
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_OFFSET 16'hbf4
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_FLD_VAL 4:0
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CPLX_BURST_ARRAY22_WIDTH 5

/* PRBS_MAX_ROW_COL */
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_OFFSET 16'hbf8
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_MAX_ROW 17:0
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_MAX_ROW_WIDTH 18
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_MAX_COL 24:18
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_MAX_COL_WIDTH 7
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_RESERVED 31:25
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_FLD_RESERVED_WIDTH 7
`define DDRMC5_MAIN_PRBS_MAX_ROW_COL_WIDTH 25

/* PRBS_MAX_LOOPS */
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_OFFSET 16'hbfc
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_FLD_CNT 11:0
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_FLD_CNT_WIDTH 12
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_FLD_RESERVED 31:12
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_FLD_RESERVED_WIDTH 20
`define DDRMC5_MAIN_PRBS_MAX_LOOPS_WIDTH 12

/* PRBS_TREF */
`define DDRMC5_MAIN_PRBS_TREF_OFFSET 16'hc00
`define DDRMC5_MAIN_PRBS_TREF_FLD_TRFC_AB 11:0
`define DDRMC5_MAIN_PRBS_TREF_FLD_TRFC_AB_WIDTH 12
`define DDRMC5_MAIN_PRBS_TREF_FLD_TRFC_SB_PB 23:12
`define DDRMC5_MAIN_PRBS_TREF_FLD_TRFC_SB_PB_WIDTH 12
`define DDRMC5_MAIN_PRBS_TREF_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PRBS_TREF_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PRBS_TREF_WIDTH 24

/* XPI_ADDR_CFG */
`define DDRMC5_MAIN_XPI_ADDR_CFG_OFFSET 16'hc04
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_ADD_PAR_ERR_CFG 1:0
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_ADD_PAR_ERR_CFG_WIDTH 2
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_PAR_EN 2
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_PAR_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_RCD_PAR_PAT_EN 3
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_RCD_PAR_PAT_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_DDR5_2N 4
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_DDR5_2N_WIDTH 1
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_RESERVED 31:5
`define DDRMC5_MAIN_XPI_ADDR_CFG_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_XPI_ADDR_CFG_WIDTH 5

/* PHY_RDEN0 */
`define DDRMC5_MAIN_PHY_RDEN0_OFFSET 16'hc08
`define DDRMC5_MAIN_PHY_RDEN0_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN0_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN0_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN0_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN0_WIDTH 8

/* PHY_RDEN1 */
`define DDRMC5_MAIN_PHY_RDEN1_OFFSET 16'hc0c
`define DDRMC5_MAIN_PHY_RDEN1_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN1_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN1_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN1_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN1_WIDTH 8

/* PHY_RDEN2 */
`define DDRMC5_MAIN_PHY_RDEN2_OFFSET 16'hc10
`define DDRMC5_MAIN_PHY_RDEN2_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN2_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN2_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN2_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN2_WIDTH 8

/* PHY_RDEN3 */
`define DDRMC5_MAIN_PHY_RDEN3_OFFSET 16'hc14
`define DDRMC5_MAIN_PHY_RDEN3_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN3_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN3_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN3_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN3_WIDTH 8

/* PHY_RDEN4 */
`define DDRMC5_MAIN_PHY_RDEN4_OFFSET 16'hc18
`define DDRMC5_MAIN_PHY_RDEN4_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN4_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN4_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN4_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN4_WIDTH 8

/* PHY_RDEN5 */
`define DDRMC5_MAIN_PHY_RDEN5_OFFSET 16'hc1c
`define DDRMC5_MAIN_PHY_RDEN5_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN5_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN5_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN5_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN5_WIDTH 8

/* PHY_RDEN6 */
`define DDRMC5_MAIN_PHY_RDEN6_OFFSET 16'hc20
`define DDRMC5_MAIN_PHY_RDEN6_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN6_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN6_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN6_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN6_WIDTH 8

/* PHY_RDEN7 */
`define DDRMC5_MAIN_PHY_RDEN7_OFFSET 16'hc24
`define DDRMC5_MAIN_PHY_RDEN7_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN7_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN7_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN7_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN7_WIDTH 8

/* PHY_RDEN8 */
`define DDRMC5_MAIN_PHY_RDEN8_OFFSET 16'hc28
`define DDRMC5_MAIN_PHY_RDEN8_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN8_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN8_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN8_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN8_WIDTH 8

/* PHY_RDEN9 */
`define DDRMC5_MAIN_PHY_RDEN9_OFFSET 16'hc2c
`define DDRMC5_MAIN_PHY_RDEN9_FLD_DLY 7:0
`define DDRMC5_MAIN_PHY_RDEN9_FLD_DLY_WIDTH 8
`define DDRMC5_MAIN_PHY_RDEN9_FLD_RESERVED 31:8
`define DDRMC5_MAIN_PHY_RDEN9_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_PHY_RDEN9_WIDTH 8

/* READ_DATA_EARLY_ID */
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_OFFSET 16'hc30
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_FLD_OFFSET 2:0
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_FLD_OFFSET_WIDTH 3
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_FLD_RESERVED 31:3
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_READ_DATA_EARLY_ID_WIDTH 3

/* FIFO_RDEN */
`define DDRMC5_MAIN_FIFO_RDEN_OFFSET 16'hc34
`define DDRMC5_MAIN_FIFO_RDEN_FLD_DLY 6:0
`define DDRMC5_MAIN_FIFO_RDEN_FLD_DLY_WIDTH 7
`define DDRMC5_MAIN_FIFO_RDEN_FLD_RESERVED 31:7
`define DDRMC5_MAIN_FIFO_RDEN_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_FIFO_RDEN_WIDTH 7

/* PHY_RANK_READ_OVERRIDE */
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_OFFSET 16'hc38
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_STATIC_ENABLE 0
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_STATIC_ENABLE_WIDTH 1
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_STATIC_ENABLE 1
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_STATIC_ENABLE_WIDTH 1
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK0 3:2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK0_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK1 5:4
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK1_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK2 7:6
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK2_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK3 9:8
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH0_RANK3_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK0 11:10
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK0_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK1 13:12
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK1_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK2 15:14
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK2_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK3 17:16
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_CH1_RANK3_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_RESERVED 31:18
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_PHY_RANK_READ_OVERRIDE_WIDTH 18

/* XPI_READ_OFFSET */
`define DDRMC5_MAIN_XPI_READ_OFFSET_OFFSET 16'hc3c
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_PHY_RDEN 3:0
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_PHY_RDEN_WIDTH 4
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RD_RETURN_RPTR 6:4
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RD_RETURN_RPTR_WIDTH 3
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RAW_RETURN_RPTR 9:7
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RAW_RETURN_RPTR_WIDTH 3
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RMW_BP_RETURN_RPTR 12:10
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RMW_BP_RETURN_RPTR_WIDTH 3
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RDCS_EARLY 14:13
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RDCS_EARLY_WIDTH 2
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RESERVED 31:15
`define DDRMC5_MAIN_XPI_READ_OFFSET_FLD_RESERVED_WIDTH 17
`define DDRMC5_MAIN_XPI_READ_OFFSET_WIDTH 15

/* XPI_READ_DBI */
`define DDRMC5_MAIN_XPI_READ_DBI_OFFSET 16'hc40
`define DDRMC5_MAIN_XPI_READ_DBI_FLD_EN 0
`define DDRMC5_MAIN_XPI_READ_DBI_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_READ_DBI_FLD_RESERVED 31:1
`define DDRMC5_MAIN_XPI_READ_DBI_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_XPI_READ_DBI_WIDTH 1

/* XPI_IBUF_DIS_OR_HS_RX_DIS */
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_OFFSET 16'hc44
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_ENABLE 0
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_ENABLE_WIDTH 1
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_EXTEND_CNT 6:1
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_EXTEND_CNT_WIDTH 6
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_RESERVED 31:7
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_XPI_IBUF_DIS_OR_HS_RX_DIS_WIDTH 7

/* XPI_READ_NIB_ENABLE */
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_OFFSET 16'hc48
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_FLD_SEL 9:0
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_FLD_SEL_WIDTH 10
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_XPI_READ_NIB_ENABLE_WIDTH 10

/* DDR5_READ_LFSR_CFG */
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_OFFSET 16'hc4c
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_RESTART 0
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_RESTART_WIDTH 1
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_LFSR0_SEED 8:1
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_LFSR0_SEED_WIDTH 8
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_LFSR1_SEED 16:9
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_LFSR1_SEED_WIDTH 8
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DDR5_READ_LFSR_CFG_WIDTH 17

/* DDR5_READ_LFSR_INVERT_31_0 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_31_0_OFFSET 16'hc50
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_31_0_FLD_EN 31:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_31_0_FLD_EN_WIDTH 32
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_31_0_WIDTH 32

/* DDR5_READ_LFSR_INVERT_39_32 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_OFFSET 16'hc54
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_FLD_EN 7:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_FLD_EN_WIDTH 8
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_DDR5_READ_LFSR_INVERT_39_32_WIDTH 8

/* DDR5_READ_LFSR_OPT_31_0 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_31_0_OFFSET 16'hc58
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_31_0_FLD_OPT 31:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_31_0_FLD_OPT_WIDTH 32
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_31_0_WIDTH 32

/* DDR5_READ_LFSR_OPT_39_32 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_OFFSET 16'hc5c
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_FLD_OPT 7:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_FLD_OPT_WIDTH 8
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_DDR5_READ_LFSR_OPT_39_32_WIDTH 8

/* DDR5_READ_LFSR_PAT_31_0 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_31_0_OFFSET 16'hc60
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_31_0_FLD_PAT 31:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_31_0_FLD_PAT_WIDTH 32
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_31_0_WIDTH 32

/* DDR5_READ_LFSR_PAT_39_32 */
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_OFFSET 16'hc64
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_FLD_PAT 7:0
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_FLD_PAT_WIDTH 8
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_DDR5_READ_LFSR_PAT_39_32_WIDTH 8

/* DDR5_SPARE_DYN_CFG0 */
`define DDRMC5_MAIN_DDR5_SPARE_DYN_CFG0_OFFSET 16'hc68
`define DDRMC5_MAIN_DDR5_SPARE_DYN_CFG0_FLD_SPARE 31:0
`define DDRMC5_MAIN_DDR5_SPARE_DYN_CFG0_FLD_SPARE_WIDTH 32
`define DDRMC5_MAIN_DDR5_SPARE_DYN_CFG0_WIDTH 32

/* REG_COM_0 */
`define DDRMC5_MAIN_REG_COM_0_OFFSET 16'hc6c
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_REQ 0
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_REQ_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_ACK 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_ACK_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_DONE 2
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_DONE_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_ERROR 3
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_ENTER_ERROR_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_REQ 4
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_REQ_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_ACK 5
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_ACK_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_DONE 6
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_DONE_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_ERROR 7
`define DDRMC5_MAIN_REG_COM_0_FLD_SELF_REFRESH_EXIT_ERROR_WIDTH 1
`define DDRMC5_MAIN_REG_COM_0_FLD_RESERVED 31:8
`define DDRMC5_MAIN_REG_COM_0_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_REG_COM_0_WIDTH 8

/* REG_COM_4 */
`define DDRMC5_MAIN_REG_COM_4_OFFSET 16'hc70
`define DDRMC5_MAIN_REG_COM_4_FLD_DRAM_MODE_REPORT 4:0
`define DDRMC5_MAIN_REG_COM_4_FLD_DRAM_MODE_REPORT_WIDTH 5
`define DDRMC5_MAIN_REG_COM_4_FLD_RESERVED 31:5
`define DDRMC5_MAIN_REG_COM_4_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_REG_COM_4_WIDTH 5

/* REG_COM_5 */
`define DDRMC5_MAIN_REG_COM_5_OFFSET 16'hc74
`define DDRMC5_MAIN_REG_COM_5_FLD_ENABLE_CRYPTO_MEM_FILL 0
`define DDRMC5_MAIN_REG_COM_5_FLD_ENABLE_CRYPTO_MEM_FILL_WIDTH 1
`define DDRMC5_MAIN_REG_COM_5_FLD_CRYPTO_FILL_EN 1
`define DDRMC5_MAIN_REG_COM_5_FLD_CRYPTO_FILL_EN_WIDTH 1
`define DDRMC5_MAIN_REG_COM_5_FLD_CRYPTO_FILL_DONE 2
`define DDRMC5_MAIN_REG_COM_5_FLD_CRYPTO_FILL_DONE_WIDTH 1
`define DDRMC5_MAIN_REG_COM_5_FLD_DDRMC_BUSY 3
`define DDRMC5_MAIN_REG_COM_5_FLD_DDRMC_BUSY_WIDTH 1
`define DDRMC5_MAIN_REG_COM_5_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_COM_5_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_COM_5_WIDTH 4

/* REG_MRS_3 */
`define DDRMC5_MAIN_REG_MRS_3_OFFSET 16'hc78
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_MRA_DDR5 7:0
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_MRA_DDR5_WIDTH 8
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_OPCODE 15:8
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_OPCODE_WIDTH 8
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_MA_LPDDR5 21:16
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_CMD_MA_LPDDR5_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_PREA_SKIP_DDR5 22
`define DDRMC5_MAIN_REG_MRS_3_FLD_MR_PREA_SKIP_DDR5_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_3_FLD_RESERVED 31:23
`define DDRMC5_MAIN_REG_MRS_3_FLD_RESERVED_WIDTH 9
`define DDRMC5_MAIN_REG_MRS_3_WIDTH 23

/* REG_MRS_4 */
`define DDRMC5_MAIN_REG_MRS_4_OFFSET 16'hc7c
`define DDRMC5_MAIN_REG_MRS_4_FLD_MR_CMD_TYPE 2:0
`define DDRMC5_MAIN_REG_MRS_4_FLD_MR_CMD_TYPE_WIDTH 3
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_ADDR 8:3
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_ADDR_WIDTH 6
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_CS 12:9
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_CS_WIDTH 4
`define DDRMC5_MAIN_REG_MRS_4_FLD_RESERVED 14:13
`define DDRMC5_MAIN_REG_MRS_4_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_MIRROR 15
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_MIRROR_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_INVERT 16
`define DDRMC5_MAIN_REG_MRS_4_FLD_MRS_INVERT_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_4_FLD_RESERVED_1 31:17
`define DDRMC5_MAIN_REG_MRS_4_FLD_RESERVED_1_WIDTH 15
`define DDRMC5_MAIN_REG_MRS_4_WIDTH 17

/* REG_MRS_5 */
`define DDRMC5_MAIN_REG_MRS_5_OFFSET 16'hc80
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_START_0 0
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_START_0_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_BUSY_0 1
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_BUSY_0_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_DONE_0 2
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_DONE_0_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_ERROR_0 3
`define DDRMC5_MAIN_REG_MRS_5_FLD_MRS_COMMAND_ERROR_0_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_5_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_MRS_5_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_MRS_5_WIDTH 4

/* REG_MRS_6 */
`define DDRMC5_MAIN_REG_MRS_6_OFFSET 16'hc84
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_START_1 0
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_START_1_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_BUSY_1 1
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_BUSY_1_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_DONE_1 2
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_DONE_1_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_ERROR_1 3
`define DDRMC5_MAIN_REG_MRS_6_FLD_MRS_COMMAND_ERROR_1_WIDTH 1
`define DDRMC5_MAIN_REG_MRS_6_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_MRS_6_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_MRS_6_WIDTH 4

/* REG_SCRUB_STATUS_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_OFFSET 16'hc88
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_START 0
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_START_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_STOP 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_STOP_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_BUSY 2
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_BUSY_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_DONE 3
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_SCRUB_DONE_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH0_WIDTH 4

/* REG_SCRUB_STATUS_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_OFFSET 16'hc8c
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_START 0
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_START_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_STOP 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_STOP_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_BUSY 2
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_BUSY_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_DONE 3
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_SCRUB_DONE_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_RESERVED 31:4
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_REG_SCRUB_STATUS_CH1_WIDTH 4

/* REG_SCRUB_ADDR_LO_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH0_OFFSET 16'hc90
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH0_FLD_SCRUB_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH0_FLD_SCRUB_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH0_WIDTH 32

/* REG_SCRUB_ADDR_HI_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_OFFSET 16'hc94
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_FLD_SCRUB_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_FLD_SCRUB_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH0_WIDTH 16

/* REG_SCRUB_ADDR_LO_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH1_OFFSET 16'hc98
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH1_FLD_SCRUB_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH1_FLD_SCRUB_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_ADDR_LO_CH1_WIDTH 32

/* REG_SCRUB_ADDR_HI_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_OFFSET 16'hc9c
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_FLD_SCRUB_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_FLD_SCRUB_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_ADDR_HI_CH1_WIDTH 16

/* REG_SCRUB_LOOP_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_OFFSET 16'hca0
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_FLD_NUM_FULL_SCRUB 7:0
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_FLD_NUM_FULL_SCRUB_WIDTH 8
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_FLD_RESERVED 31:8
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH0_WIDTH 8

/* REG_SCRUB_LOOP_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_OFFSET 16'hca4
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_FLD_NUM_FULL_SCRUB 7:0
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_FLD_NUM_FULL_SCRUB_WIDTH 8
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_FLD_RESERVED 31:8
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_REG_SCRUB_LOOP_CH1_WIDTH 8

/* REG_SCRUB_EVENT_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_OFFSET 16'hca8
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_SCRUB_TO_EVENT 0
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_SCRUB_TO_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_PER_RD_TO_EVENT 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_PER_RD_TO_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_ASYNC_FIFO_FULL 2
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_ASYNC_FIFO_FULL_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_TXN_COUNTER_ROLLOVER 3
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_TXN_COUNTER_ROLLOVER_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_MISSED_SCRUB_EVENT 4
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_MISSED_SCRUB_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_MISSED_PER_RD_EVENT 5
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_MISSED_PER_RD_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_RESERVED 31:6
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_FLD_RESERVED_WIDTH 26
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH0_WIDTH 6

/* REG_SCRUB_EVENT_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_OFFSET 16'hcac
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_SCRUB_TO_EVENT 0
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_SCRUB_TO_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_PER_RD_TO_EVENT 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_PER_RD_TO_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_ASYNC_FIFO_FULL 2
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_ASYNC_FIFO_FULL_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_TXN_COUNTER_ROLLOVER 3
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_TXN_COUNTER_ROLLOVER_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_MISSED_SCRUB_EVENT 4
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_MISSED_SCRUB_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_MISSED_PER_RD_EVENT 5
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_MISSED_PER_RD_EVENT_WIDTH 1
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_RESERVED 31:6
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_FLD_RESERVED_WIDTH 26
`define DDRMC5_MAIN_REG_SCRUB_EVENT_CH1_WIDTH 6

/* REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH0_OFFSET 16'hcb0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH0_FLD_MISSED_SCRUB_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH0_FLD_MISSED_SCRUB_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH0_WIDTH 32

/* REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_OFFSET 16'hcb4
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_FLD_MISSED_SCRUB_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_FLD_MISSED_SCRUB_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH0_WIDTH 16

/* REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH1_OFFSET 16'hcb8
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH1_FLD_MISSED_SCRUB_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH1_FLD_MISSED_SCRUB_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_LO_CH1_WIDTH 32

/* REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_OFFSET 16'hcbc
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_FLD_MISSED_SCRUB_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_FLD_MISSED_SCRUB_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_ADDR_HI_CH1_WIDTH 16

/* REG_SCRUB_MISSED_SCRUB_PARA_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH0_OFFSET 16'hcc0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH0_FLD_MISSED_SCRUB_PARAMETER 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH0_FLD_MISSED_SCRUB_PARAMETER_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH0_WIDTH 32

/* REG_SCRUB_MISSED_SCRUB_PARA_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH1_OFFSET 16'hcc4
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH1_FLD_MISSED_SCRUB_PARAMETER 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH1_FLD_MISSED_SCRUB_PARAMETER_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_SCRUB_PARA_CH1_WIDTH 32

/* REG_SCRUB_MISSED_PER_RD_LO_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH0_OFFSET 16'hcc8
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH0_FLD_MISSED_PER_RD_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH0_FLD_MISSED_PER_RD_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH0_WIDTH 32

/* REG_SCRUB_MISSED_PER_RD_HI_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_OFFSET 16'hccc
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_FLD_MISSED_PER_RD_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_FLD_MISSED_PER_RD_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH0_WIDTH 16

/* REG_SCRUB_MISSED_PER_RD_LO_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH1_OFFSET 16'hcd0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH1_FLD_MISSED_PER_RD_CURRENT_OFFSET 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH1_FLD_MISSED_PER_RD_CURRENT_OFFSET_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_LO_CH1_WIDTH 32

/* REG_SCRUB_MISSED_PER_RD_HI_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_OFFSET 16'hcd4
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_FLD_MISSED_PER_RD_CURRENT_OFFSET 15:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_FLD_MISSED_PER_RD_CURRENT_OFFSET_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_HI_CH1_WIDTH 16

/* REG_SCRUB_MISSED_PER_RD_PARA_CH0 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH0_OFFSET 16'hcd8
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH0_FLD_MISSED_PER_RD_PARAMETER 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH0_FLD_MISSED_PER_RD_PARAMETER_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH0_WIDTH 32

/* REG_SCRUB_MISSED_PER_RD_PARA_CH1 */
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH1_OFFSET 16'hcdc
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH1_FLD_MISSED_PER_RD_PARAMETER 31:0
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH1_FLD_MISSED_PER_RD_PARAMETER_WIDTH 32
`define DDRMC5_MAIN_REG_SCRUB_MISSED_PER_RD_PARA_CH1_WIDTH 32

/* DC_QUEUE_STATUS */
`define DDRMC5_MAIN_DC_QUEUE_STATUS_OFFSET 16'hce0
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL0 0
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL0_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL0_STKY 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL0_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY0 2
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY0_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY0_STKY 3
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY0_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_SKIP0_STKY 4
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_SKIP0_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_STARVED0_STKY 5
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_STARVED0_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_RESERVED 15:6
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_RESERVED_WIDTH 10
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL1 16
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL1_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL1_STKY 17
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_FULL1_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY1 18
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY1_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY1_STKY 19
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_EMPTY1_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_SKIP1_STKY 20
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_SKIP1_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_STARVED1_STKY 21
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_STARVED1_STKY_WIDTH 1
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_RESERVED_1 31:22
`define DDRMC5_MAIN_DC_QUEUE_STATUS_FLD_RESERVED_1_WIDTH 10
`define DDRMC5_MAIN_DC_QUEUE_STATUS_WIDTH 22

/* WRCS_STARTUP_NIB_DONE */
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_OFFSET 16'hce4
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_CH0 9:0
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_CH0_WIDTH 10
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_CH1 19:10
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_CH1_WIDTH 10
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_RESERVED 31:20
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_WRCS_STARTUP_NIB_DONE_WIDTH 20

/* PHY_OE_NIB_ERR */
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_OFFSET 16'hce8
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH0_DLY_UNDERFLOW 9:0
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH0_DLY_UNDERFLOW_WIDTH 10
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH1_DLY_UNDERFLOW 19:10
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH1_DLY_UNDERFLOW_WIDTH 10
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH0_DLY_OVERFLOW 29:20
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH0_DLY_OVERFLOW_WIDTH 10
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH1_DLY_OVERFLOW 30
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_CH1_DLY_OVERFLOW_WIDTH 1
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_RESERVED 31
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_PHY_OE_NIB_ERR_WIDTH 31

/* PHY_WDATA_ERR */
`define DDRMC5_MAIN_PHY_WDATA_ERR_OFFSET 16'hcec
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_CH0_DLY_UNDERFLOW 0
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_CH0_DLY_UNDERFLOW_WIDTH 1
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_CH1_DLY_UNDERFLOW 1
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_CH1_DLY_UNDERFLOW_WIDTH 1
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_RESERVED 31:2
`define DDRMC5_MAIN_PHY_WDATA_ERR_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_PHY_WDATA_ERR_WIDTH 2

/* XPI_DYN_RANK */
`define DDRMC5_MAIN_XPI_DYN_RANK_OFFSET 16'hcf0
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_BUSY 0
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_BUSY_WIDTH 1
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_DONE_CNT 2:1
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_DONE_CNT_WIDTH 2
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_DBG 4:3
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH0_DBG_WIDTH 2
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_BUSY 5
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_BUSY_WIDTH 1
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_DONE_CNT 7:6
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_DONE_CNT_WIDTH 2
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_DBG 9:8
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_CH1_DBG_WIDTH 2
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_RESERVED 31:10
`define DDRMC5_MAIN_XPI_DYN_RANK_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_XPI_DYN_RANK_WIDTH 10

/* PHY_OE_NIB0 */
`define DDRMC5_MAIN_PHY_OE_NIB0_OFFSET 16'hcf4
`define DDRMC5_MAIN_PHY_OE_NIB0_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB0_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB0_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB0_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB0_WIDTH 3

/* PHY_OE_NIB1 */
`define DDRMC5_MAIN_PHY_OE_NIB1_OFFSET 16'hcf8
`define DDRMC5_MAIN_PHY_OE_NIB1_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB1_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB1_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB1_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB1_WIDTH 3

/* PHY_OE_NIB2 */
`define DDRMC5_MAIN_PHY_OE_NIB2_OFFSET 16'hcfc
`define DDRMC5_MAIN_PHY_OE_NIB2_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB2_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB2_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB2_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB2_WIDTH 3

/* PHY_OE_NIB3 */
`define DDRMC5_MAIN_PHY_OE_NIB3_OFFSET 16'hd00
`define DDRMC5_MAIN_PHY_OE_NIB3_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB3_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB3_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB3_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB3_WIDTH 3

/* PHY_OE_NIB4 */
`define DDRMC5_MAIN_PHY_OE_NIB4_OFFSET 16'hd04
`define DDRMC5_MAIN_PHY_OE_NIB4_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB4_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB4_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB4_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB4_WIDTH 3

/* PHY_OE_NIB5 */
`define DDRMC5_MAIN_PHY_OE_NIB5_OFFSET 16'hd08
`define DDRMC5_MAIN_PHY_OE_NIB5_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB5_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB5_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB5_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB5_WIDTH 3

/* PHY_OE_NIB6 */
`define DDRMC5_MAIN_PHY_OE_NIB6_OFFSET 16'hd0c
`define DDRMC5_MAIN_PHY_OE_NIB6_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB6_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB6_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB6_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB6_WIDTH 3

/* PHY_OE_NIB7 */
`define DDRMC5_MAIN_PHY_OE_NIB7_OFFSET 16'hd10
`define DDRMC5_MAIN_PHY_OE_NIB7_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB7_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB7_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB7_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB7_WIDTH 3

/* PHY_OE_NIB8 */
`define DDRMC5_MAIN_PHY_OE_NIB8_OFFSET 16'hd14
`define DDRMC5_MAIN_PHY_OE_NIB8_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB8_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB8_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB8_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB8_WIDTH 3

/* PHY_OE_NIB9 */
`define DDRMC5_MAIN_PHY_OE_NIB9_OFFSET 16'hd18
`define DDRMC5_MAIN_PHY_OE_NIB9_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_OE_NIB9_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_OE_NIB9_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_OE_NIB9_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_OE_NIB9_WIDTH 3

/* CAL_STATUS */
`define DDRMC5_MAIN_CAL_STATUS_OFFSET 16'hd1c
`define DDRMC5_MAIN_CAL_STATUS_FLD_INIT_DONE 0
`define DDRMC5_MAIN_CAL_STATUS_FLD_INIT_DONE_WIDTH 1
`define DDRMC5_MAIN_CAL_STATUS_FLD_CAL_DONE 1
`define DDRMC5_MAIN_CAL_STATUS_FLD_CAL_DONE_WIDTH 1
`define DDRMC5_MAIN_CAL_STATUS_FLD_RESERVED 31:2
`define DDRMC5_MAIN_CAL_STATUS_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_CAL_STATUS_WIDTH 2

/* BL8_NIBBLE0 */
`define DDRMC5_MAIN_BL8_NIBBLE0_OFFSET 16'hd20
`define DDRMC5_MAIN_BL8_NIBBLE0_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE0_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE0_WIDTH 32

/* BL8_NIBBLE1 */
`define DDRMC5_MAIN_BL8_NIBBLE1_OFFSET 16'hd24
`define DDRMC5_MAIN_BL8_NIBBLE1_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE1_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE1_WIDTH 32

/* BL8_NIBBLE2 */
`define DDRMC5_MAIN_BL8_NIBBLE2_OFFSET 16'hd28
`define DDRMC5_MAIN_BL8_NIBBLE2_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE2_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE2_WIDTH 32

/* BL8_NIBBLE3 */
`define DDRMC5_MAIN_BL8_NIBBLE3_OFFSET 16'hd2c
`define DDRMC5_MAIN_BL8_NIBBLE3_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE3_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE3_WIDTH 32

/* BL8_NIBBLE4 */
`define DDRMC5_MAIN_BL8_NIBBLE4_OFFSET 16'hd30
`define DDRMC5_MAIN_BL8_NIBBLE4_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE4_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE4_WIDTH 32

/* BL8_NIBBLE5 */
`define DDRMC5_MAIN_BL8_NIBBLE5_OFFSET 16'hd34
`define DDRMC5_MAIN_BL8_NIBBLE5_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE5_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE5_WIDTH 32

/* BL8_NIBBLE6 */
`define DDRMC5_MAIN_BL8_NIBBLE6_OFFSET 16'hd38
`define DDRMC5_MAIN_BL8_NIBBLE6_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE6_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE6_WIDTH 32

/* BL8_NIBBLE7 */
`define DDRMC5_MAIN_BL8_NIBBLE7_OFFSET 16'hd3c
`define DDRMC5_MAIN_BL8_NIBBLE7_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE7_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE7_WIDTH 32

/* BL8_NIBBLE8 */
`define DDRMC5_MAIN_BL8_NIBBLE8_OFFSET 16'hd40
`define DDRMC5_MAIN_BL8_NIBBLE8_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE8_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE8_WIDTH 32

/* BL8_NIBBLE9 */
`define DDRMC5_MAIN_BL8_NIBBLE9_OFFSET 16'hd44
`define DDRMC5_MAIN_BL8_NIBBLE9_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL8_NIBBLE9_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL8_NIBBLE9_WIDTH 32

/* COMPARE_CLEAR */
`define DDRMC5_MAIN_COMPARE_CLEAR_OFFSET 16'hd48
`define DDRMC5_MAIN_COMPARE_CLEAR_FLD_VAL 0
`define DDRMC5_MAIN_COMPARE_CLEAR_FLD_VAL_WIDTH 1
`define DDRMC5_MAIN_COMPARE_CLEAR_FLD_RESERVED 31:1
`define DDRMC5_MAIN_COMPARE_CLEAR_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_COMPARE_CLEAR_WIDTH 1

/* COMPARE_CONFIG */
`define DDRMC5_MAIN_COMPARE_CONFIG_OFFSET 16'hd4c
`define DDRMC5_MAIN_COMPARE_CONFIG_FLD_ERR_EN 0
`define DDRMC5_MAIN_COMPARE_CONFIG_FLD_ERR_EN_WIDTH 1
`define DDRMC5_MAIN_COMPARE_CONFIG_FLD_RESERVED 31:1
`define DDRMC5_MAIN_COMPARE_CONFIG_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_COMPARE_CONFIG_WIDTH 1

/* ERR_PER_BIT_ANY_REDGE_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_31_0_OFFSET 16'hd50
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_31_0_WIDTH 32

/* ERR_PER_BIT_ANY_REDGE_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_OFFSET 16'hd54
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_39_32_WIDTH 8

/* ERR_PER_BIT_ALL_REDGES_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_31_0_OFFSET 16'hd58
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_31_0_WIDTH 32

/* ERR_PER_BIT_ALL_REDGES_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_OFFSET 16'hd5c
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_REDGES_39_32_WIDTH 8

/* ERR_PER_BIT_ANY_FEDGE_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_31_0_OFFSET 16'hd60
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_31_0_WIDTH 32

/* ERR_PER_BIT_ANY_FEDGE_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_OFFSET 16'hd64
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_FEDGE_39_32_WIDTH 8

/* ERR_PER_BIT_ALL_FEDGES_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_31_0_OFFSET 16'hd68
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_31_0_WIDTH 32

/* ERR_PER_BIT_ALL_FEDGES_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_OFFSET 16'hd6c
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_FEDGES_39_32_WIDTH 8

/* ERR_PER_BIT_ANY_EDGE_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_OFFSET 16'hd70
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_WIDTH 32

/* ERR_PER_BIT_ANY_EDGE_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_OFFSET 16'hd74
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_WIDTH 8

/* ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_31_0_OFFSET 16'hd78
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_31_0_WIDTH 32

/* ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_OFFSET 16'hd7c
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_REDGE_AND_ANY_FEDGE_39_32_WIDTH 8

/* ERR_PER_BIT_ALL_EDGES_31_0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_31_0_OFFSET 16'hd80
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_31_0_WIDTH 32

/* ERR_PER_BIT_ALL_EDGES_39_32 */
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_OFFSET 16'hd84
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ALL_EDGES_39_32_WIDTH 8

/* ERR_PER_NIB_ANY_BIT_ANY_REDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_OFFSET 16'hd88
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_REDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ANY_REDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_OFFSET 16'hd8c
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_REDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ALL_REDGES */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_OFFSET 16'hd90
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_REDGES_WIDTH 10

/* ERR_PER_NIB_ANY_BIT_ANY_FEDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_OFFSET 16'hd94
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_FEDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ANY_FEDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_OFFSET 16'hd98
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_FEDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ALL_FEDGES */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_OFFSET 16'hd9c
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_FEDGES_WIDTH 10

/* ERR_PER_NIB_ANY_BIT_ANY_EDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_OFFSET 16'hda0
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ANY_BIT_ANY_EDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ANY_EDGE */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_OFFSET 16'hda4
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ANY_EDGE_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_BOTH_EDGES */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_OFFSET 16'hda8
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_BOTH_EDGES_WIDTH 10

/* ERR_PER_NIB_ALL_BITS_ALL_EDGES */
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_OFFSET 16'hdac
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_FLD_VAL 9:0
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_FLD_VAL_WIDTH 10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_FLD_RESERVED 31:10
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_ERR_PER_NIB_ALL_BITS_ALL_EDGES_WIDTH 10

/* ERR_PER_BYT_ANY_BIT_ANY_REDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_OFFSET 16'hdb0
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_REDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ANY_REDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_OFFSET 16'hdb4
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_REDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ALL_REDGES */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_OFFSET 16'hdb8
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_REDGES_WIDTH 5

/* ERR_PER_BYT_ANY_BIT_ANY_FEDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_OFFSET 16'hdbc
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_FEDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ANY_FEDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_OFFSET 16'hdc0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_FEDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ALL_FEDGES */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_OFFSET 16'hdc4
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_FEDGES_WIDTH 5

/* ERR_PER_BYT_ANY_BIT_ANY_EDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_OFFSET 16'hdc8
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ANY_BIT_ANY_EDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ANY_EDGE */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_OFFSET 16'hdcc
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ANY_EDGE_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_BOTH_EDGES */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_OFFSET 16'hdd0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_BOTH_EDGES_WIDTH 5

/* ERR_PER_BYT_ALL_BITS_ALL_EDGES */
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_OFFSET 16'hdd4
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_FLD_VAL 4:0
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_FLD_RESERVED 31:5
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_ERR_PER_BYT_ALL_BITS_ALL_EDGES_WIDTH 5

/* COMPARE_DATA_STABLE_NIBBLE */
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_OFFSET 16'hdd8
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_FLD_VAL 19:0
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_FLD_VAL_WIDTH 20
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_FLD_RESERVED 31:20
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_COMPARE_DATA_STABLE_NIBBLE_WIDTH 20

/* COMPARE_CA_SAMPLE_STATUS_COMP0 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_OFFSET 16'hddc
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP0_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP1 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_OFFSET 16'hde0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP1_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP2 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_OFFSET 16'hde4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP2_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP3 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_OFFSET 16'hde8
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP3_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP4 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_OFFSET 16'hdec
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP4_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP5 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_OFFSET 16'hdf0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP5_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP6 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_OFFSET 16'hdf4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP6_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP7 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_OFFSET 16'hdf8
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP7_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP8 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_OFFSET 16'hdfc
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP8_WIDTH 28

/* COMPARE_CA_SAMPLE_STATUS_COMP9 */
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_OFFSET 16'he00
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_STABLE0 13:0
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_STABLE0_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_STABLE1 27:14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_STABLE1_WIDTH 14
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_RESERVED 31:28
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_FLD_RESERVED_WIDTH 4
`define DDRMC5_MAIN_COMPARE_CA_SAMPLE_STATUS_COMP9_WIDTH 28

/* ERR_PER_BIT_ANY_EDGE_31_0_DQ0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_DQ0_OFFSET 16'he04
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_DQ0_FLD_VAL 31:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_DQ0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_31_0_DQ0_WIDTH 32

/* ERR_PER_BIT_ANY_EDGE_39_32_DQ0 */
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_OFFSET 16'he08
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_FLD_VAL 7:0
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_FLD_VAL_WIDTH 8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ERR_PER_BIT_ANY_EDGE_39_32_DQ0_WIDTH 8

/* ERR_PER_BEAT_CMPR_MASK_BL16 */
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_OFFSET 16'he0c
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_BEATS 15:0
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_BEATS_WIDTH 16
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_CMP_TYPE 16
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_CMP_TYPE_WIDTH 1
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_RESERVED 31:17
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_ERR_PER_BEAT_CMPR_MASK_BL16_WIDTH 17

/* CMD2CMPR_DLY */
`define DDRMC5_MAIN_CMD2CMPR_DLY_OFFSET 16'he10
`define DDRMC5_MAIN_CMD2CMPR_DLY_FLD_VAL 4:0
`define DDRMC5_MAIN_CMD2CMPR_DLY_FLD_VAL_WIDTH 5
`define DDRMC5_MAIN_CMD2CMPR_DLY_FLD_RESERVED 31:5
`define DDRMC5_MAIN_CMD2CMPR_DLY_FLD_RESERVED_WIDTH 27
`define DDRMC5_MAIN_CMD2CMPR_DLY_WIDTH 5

/* PHY_DATA_NIB0 */
`define DDRMC5_MAIN_PHY_DATA_NIB0_OFFSET 16'he14
`define DDRMC5_MAIN_PHY_DATA_NIB0_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB0_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB0_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB0_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB0_WIDTH 3

/* PHY_DATA_NIB1 */
`define DDRMC5_MAIN_PHY_DATA_NIB1_OFFSET 16'he18
`define DDRMC5_MAIN_PHY_DATA_NIB1_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB1_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB1_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB1_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB1_WIDTH 3

/* PHY_DATA_NIB2 */
`define DDRMC5_MAIN_PHY_DATA_NIB2_OFFSET 16'he1c
`define DDRMC5_MAIN_PHY_DATA_NIB2_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB2_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB2_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB2_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB2_WIDTH 3

/* PHY_DATA_NIB3 */
`define DDRMC5_MAIN_PHY_DATA_NIB3_OFFSET 16'he20
`define DDRMC5_MAIN_PHY_DATA_NIB3_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB3_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB3_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB3_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB3_WIDTH 3

/* PHY_DATA_NIB4 */
`define DDRMC5_MAIN_PHY_DATA_NIB4_OFFSET 16'he24
`define DDRMC5_MAIN_PHY_DATA_NIB4_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB4_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB4_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB4_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB4_WIDTH 3

/* PHY_DATA_NIB5 */
`define DDRMC5_MAIN_PHY_DATA_NIB5_OFFSET 16'he28
`define DDRMC5_MAIN_PHY_DATA_NIB5_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB5_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB5_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB5_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB5_WIDTH 3

/* PHY_DATA_NIB6 */
`define DDRMC5_MAIN_PHY_DATA_NIB6_OFFSET 16'he2c
`define DDRMC5_MAIN_PHY_DATA_NIB6_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB6_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB6_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB6_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB6_WIDTH 3

/* PHY_DATA_NIB7 */
`define DDRMC5_MAIN_PHY_DATA_NIB7_OFFSET 16'he30
`define DDRMC5_MAIN_PHY_DATA_NIB7_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB7_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB7_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB7_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB7_WIDTH 3

/* PHY_DATA_NIB8 */
`define DDRMC5_MAIN_PHY_DATA_NIB8_OFFSET 16'he34
`define DDRMC5_MAIN_PHY_DATA_NIB8_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB8_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB8_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB8_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB8_WIDTH 3

/* PHY_DATA_NIB9 */
`define DDRMC5_MAIN_PHY_DATA_NIB9_OFFSET 16'he38
`define DDRMC5_MAIN_PHY_DATA_NIB9_FLD_DLY 2:0
`define DDRMC5_MAIN_PHY_DATA_NIB9_FLD_DLY_WIDTH 3
`define DDRMC5_MAIN_PHY_DATA_NIB9_FLD_RESERVED 31:3
`define DDRMC5_MAIN_PHY_DATA_NIB9_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_PHY_DATA_NIB9_WIDTH 3

/* ECCW0_FLIP_CONTROL */
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_OFFSET 16'he3c
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_00 0
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_00_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_01 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_01_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_02 2
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_02_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_03 3
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_03_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_10 4
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_10_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_11 5
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_11_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_12 6
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_12_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_13 7
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_FLIP_ENABLE_13_WIDTH 1
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCW0_FLIP_CONTROL_WIDTH 8

/* ECCW0_FLIP0 */
`define DDRMC5_MAIN_ECCW0_FLIP0_OFFSET 16'he40
`define DDRMC5_MAIN_ECCW0_FLIP0_FLD_FLIP 31:0
`define DDRMC5_MAIN_ECCW0_FLIP0_FLD_FLIP_WIDTH 32
`define DDRMC5_MAIN_ECCW0_FLIP0_WIDTH 32

/* ECCW0_FLIP1 */
`define DDRMC5_MAIN_ECCW0_FLIP1_OFFSET 16'he44
`define DDRMC5_MAIN_ECCW0_FLIP1_FLD_FLIP 31:0
`define DDRMC5_MAIN_ECCW0_FLIP1_FLD_FLIP_WIDTH 32
`define DDRMC5_MAIN_ECCW0_FLIP1_WIDTH 32

/* ECCW0_FLIP2 */
`define DDRMC5_MAIN_ECCW0_FLIP2_OFFSET 16'he48
`define DDRMC5_MAIN_ECCW0_FLIP2_FLD_FLIP 14:0
`define DDRMC5_MAIN_ECCW0_FLIP2_FLD_FLIP_WIDTH 15
`define DDRMC5_MAIN_ECCW0_FLIP2_FLD_RESERVED 31:15
`define DDRMC5_MAIN_ECCW0_FLIP2_FLD_RESERVED_WIDTH 17
`define DDRMC5_MAIN_ECCW0_FLIP2_WIDTH 15

/* ECCW1_FLIP_CONTROL */
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_OFFSET 16'he4c
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_00 0
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_00_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_01 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_01_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_02 2
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_02_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_03 3
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_03_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_10 4
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_10_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_11 5
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_11_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_12 6
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_12_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_13 7
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_FLIP_ENABLE_13_WIDTH 1
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCW1_FLIP_CONTROL_WIDTH 8

/* ECCW1_FLIP0 */
`define DDRMC5_MAIN_ECCW1_FLIP0_OFFSET 16'he50
`define DDRMC5_MAIN_ECCW1_FLIP0_FLD_FLIP 31:0
`define DDRMC5_MAIN_ECCW1_FLIP0_FLD_FLIP_WIDTH 32
`define DDRMC5_MAIN_ECCW1_FLIP0_WIDTH 32

/* ECCW1_FLIP1 */
`define DDRMC5_MAIN_ECCW1_FLIP1_OFFSET 16'he54
`define DDRMC5_MAIN_ECCW1_FLIP1_FLD_FLIP 31:0
`define DDRMC5_MAIN_ECCW1_FLIP1_FLD_FLIP_WIDTH 32
`define DDRMC5_MAIN_ECCW1_FLIP1_WIDTH 32

/* ECCW1_FLIP2 */
`define DDRMC5_MAIN_ECCW1_FLIP2_OFFSET 16'he58
`define DDRMC5_MAIN_ECCW1_FLIP2_FLD_FLIP 14:0
`define DDRMC5_MAIN_ECCW1_FLIP2_FLD_FLIP_WIDTH 15
`define DDRMC5_MAIN_ECCW1_FLIP2_FLD_RESERVED 31:15
`define DDRMC5_MAIN_ECCW1_FLIP2_FLD_RESERVED_WIDTH 17
`define DDRMC5_MAIN_ECCW1_FLIP2_WIDTH 15

/* ECCR0_CORR_ERR_STATUS */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_OFFSET 16'he5c
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR00 0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR00_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR01 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR01_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR02 2
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR02_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR03 3
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR03_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR10 4
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR10_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR11 5
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR11_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR12 6
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR12_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR13 7
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_CORR13_WIDTH 1
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCR0_CORR_ERR_STATUS_WIDTH 8

/* ECCR0_CORR_ERR_ADD_LO */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_LO_OFFSET 16'he60
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO 31:0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO_WIDTH 32
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_LO_WIDTH 32

/* ECCR0_CORR_ERR_ADD_HI */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_OFFSET 16'he64
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI 10:0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI_WIDTH 11
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_FLD_RESERVED 31:11
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_ECCR0_CORR_ERR_ADD_HI_WIDTH 11

/* ECCR0_CORR_ERR_DATA_LO */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_LO_OFFSET 16'he68
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW 31:0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW_WIDTH 32
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_LO_WIDTH 32

/* ECCR0_CORR_ERR_DATA_HI */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_HI_OFFSET 16'he6c
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI 31:0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI_WIDTH 32
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_HI_WIDTH 32

/* ECCR0_CORR_ERR_DATA_PAR */
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_OFFSET 16'he70
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR 15:0
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR_WIDTH 16
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ECCR0_CORR_ERR_DATA_PAR_WIDTH 16

/* ECCR0_UNCORR_ERR_STATUS */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_OFFSET 16'he74
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR00 0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR00_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR01 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR01_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR02 2
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR02_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR03 3
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR03_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR10 4
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR10_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR11 5
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR11_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR12 6
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR12_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR13 7
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_UNCORR13_WIDTH 1
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_STATUS_WIDTH 8

/* ECCR0_UNCORR_ERR_ADD_LO */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_LO_OFFSET 16'he78
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO 31:0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO_WIDTH 32
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_LO_WIDTH 32

/* ECCR0_UNCORR_ERR_ADD_HI */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_OFFSET 16'he7c
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI 10:0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI_WIDTH 11
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_FLD_RESERVED 31:11
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_ADD_HI_WIDTH 11

/* ECCR0_UNCORR_ERR_DATA_LO */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_LO_OFFSET 16'he80
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW 31:0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW_WIDTH 32
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_LO_WIDTH 32

/* ECCR0_UNCORR_ERR_DATA_HI */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_HI_OFFSET 16'he84
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI 31:0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI_WIDTH 32
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_HI_WIDTH 32

/* ECCR0_UNCORR_ERR_DATA_PAR */
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_OFFSET 16'he88
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR 15:0
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR_WIDTH 16
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ECCR0_UNCORR_ERR_DATA_PAR_WIDTH 16

/* ECCR1_CORR_ERR_STATUS */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_OFFSET 16'he8c
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR00 0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR00_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR01 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR01_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR02 2
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR02_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR03 3
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR03_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR10 4
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR10_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR11 5
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR11_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR12 6
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR12_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR13 7
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_CORR13_WIDTH 1
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCR1_CORR_ERR_STATUS_WIDTH 8

/* ECCR1_CORR_ERR_ADD_LO */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_LO_OFFSET 16'he90
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO 31:0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO_WIDTH 32
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_LO_WIDTH 32

/* ECCR1_CORR_ERR_ADD_HI */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_OFFSET 16'he94
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI 10:0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI_WIDTH 11
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_FLD_RESERVED 31:11
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_ECCR1_CORR_ERR_ADD_HI_WIDTH 11

/* ECCR1_CORR_ERR_DATA_LO */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_LO_OFFSET 16'he98
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW 31:0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW_WIDTH 32
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_LO_WIDTH 32

/* ECCR1_CORR_ERR_DATA_HI */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_HI_OFFSET 16'he9c
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI 31:0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI_WIDTH 32
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_HI_WIDTH 32

/* ECCR1_CORR_ERR_DATA_PAR */
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_OFFSET 16'hea0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR 15:0
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR_WIDTH 16
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ECCR1_CORR_ERR_DATA_PAR_WIDTH 16

/* ECCR1_UNCORR_ERR_STATUS */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_OFFSET 16'hea4
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR00 0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR00_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR01 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR01_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR02 2
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR02_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR03 3
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR03_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR10 4
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR10_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR11 5
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR11_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR12 6
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR12_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR13 7
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_UNCORR13_WIDTH 1
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_STATUS_WIDTH 8

/* ECCR1_UNCORR_ERR_ADD_LO */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_LO_OFFSET 16'hea8
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO 31:0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_LO_FLD_ECC_ERR_ADD_LO_WIDTH 32
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_LO_WIDTH 32

/* ECCR1_UNCORR_ERR_ADD_HI */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_OFFSET 16'heac
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI 10:0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_FLD_ECC_ERR_ADD_HI_WIDTH 11
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_FLD_RESERVED 31:11
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_FLD_RESERVED_WIDTH 21
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_ADD_HI_WIDTH 11

/* ECCR1_UNCORR_ERR_DATA_LO */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_LO_OFFSET 16'heb0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW 31:0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_LO_FLD_ECC_ERR_DATA_LOW_WIDTH 32
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_LO_WIDTH 32

/* ECCR1_UNCORR_ERR_DATA_HI */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_HI_OFFSET 16'heb4
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI 31:0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_HI_FLD_ECC_ERR_DATA_HI_WIDTH 32
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_HI_WIDTH 32

/* ECCR1_UNCORR_ERR_DATA_PAR */
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_OFFSET 16'heb8
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR 15:0
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_FLD_ECC_ERR_DATA_PAR_WIDTH 16
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ECCR1_UNCORR_ERR_DATA_PAR_WIDTH 16

/* INTERNAL_PARITY_ERROR */
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_OFFSET 16'hebc
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_PT_PARITY_0 0
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_PT_PARITY_0_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_PT_PARITY_1 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_PT_PARITY_1_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_PARITY_0 2
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_PARITY_0_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_PARITY_1 3
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_PARITY_1_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_ACAM_PARITY_0 4
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_ACAM_PARITY_0_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_ACAM_PARITY_1 5
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_ACAM_PARITY_1_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_SAFE_TIMER_PARITY_0 6
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_SAFE_TIMER_PARITY_0_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_SAFE_TIMER_PARITY_1 7
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_SAFE_TIMER_PARITY_1_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_TIMER_PARITY_0 8
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_TIMER_PARITY_0_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_TIMER_PARITY_1 9
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_TXNQ_TIMER_PARITY_1_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_RESERVED 31:10
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_WIDTH 10

/* INTERNAL_PARITY_ERROR_INJ */
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_OFFSET 16'hec0
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_0_EN 0
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_0_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_1_EN 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_1_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_0_EN 2
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_0_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_1_EN 3
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_1_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_ACAM_PARITY_0_EN 4
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_ACAM_PARITY_0_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_ACAM_PARITY_1_EN 5
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_ACAM_PARITY_1_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_RESERVED 7:6
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_ID 15:8
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_PT_PARITY_ID_WIDTH 8
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_ID 21:16
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_TXNQ_PARITY_ID_WIDTH 6
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_RESERVED_1 31:22
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_FLD_RESERVED_1_WIDTH 10
`define DDRMC5_MAIN_INTERNAL_PARITY_ERROR_INJ_WIDTH 22

/* INTERNAL_SAFE_TIMER_PARITY_ERR_CH0 */
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_OFFSET 16'hec4
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_FLD_PARITY_ERR 19:0
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_FLD_PARITY_ERR_WIDTH 20
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_FLD_RESERVED 31:20
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH0_WIDTH 20

/* INTERNAL_SAFE_TIMER_PARITY_ERR_CH1 */
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_OFFSET 16'hec8
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_FLD_PARITY_ERR 19:0
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_FLD_PARITY_ERR_WIDTH 20
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_FLD_RESERVED 31:20
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_CH1_WIDTH 20

/* INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0 */
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_OFFSET 16'hecc
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_FLD_PARITY_ERR 16:0
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_FLD_PARITY_ERR_WIDTH 17
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_FLD_RESERVED 31:17
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH0_WIDTH 17

/* INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1 */
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_OFFSET 16'hed0
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_FLD_PARITY_ERR 16:0
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_FLD_PARITY_ERR_WIDTH 17
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_FLD_RESERVED 31:17
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_CH1_WIDTH 17

/* INTERNAL_SAFE_TIMER_PARITY_ERR_INJ */
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_OFFSET 16'hed4
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_CH1_EN 0
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_CH1_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_PARITY_EN 20:1
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_PARITY_EN_WIDTH 20
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_RESERVED 31:21
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_FLD_RESERVED_WIDTH 11
`define DDRMC5_MAIN_INTERNAL_SAFE_TIMER_PARITY_ERR_INJ_WIDTH 21

/* INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ */
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_OFFSET 16'hed8
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_CH1_EN 0
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_CH1_EN_WIDTH 1
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_PARITY_EN 17:1
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_PARITY_EN_WIDTH 17
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_RESERVED 31:18
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_INTERNAL_TXNQ_TIMER_PARITY_ERR_INJ_WIDTH 18

/* XPI_LP5_CAL */
`define DDRMC5_MAIN_XPI_LP5_CAL_OFFSET 16'hedc
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_CA_CAL_MODE_EN 0
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_CA_CAL_MODE_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_MUX_CAL_DRIVE_ADDR_CS_LIKE_DC 1
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_MUX_CAL_DRIVE_ADDR_CS_LIKE_DC_WIDTH 1
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_RESERVED 31:2
`define DDRMC5_MAIN_XPI_LP5_CAL_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_XPI_LP5_CAL_WIDTH 2

/* XPI_MAP_BITSLIP */
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_OFFSET 16'hee0
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_ADDR_EN_CH0 0
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_ADDR_EN_CH0_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_ADDR_EN_CH1 1
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_ADDR_EN_CH1_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_CS_EN_CH0 7:2
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_CS_EN_CH0_WIDTH 6
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_CS_EN_CH1 13:8
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_CS_EN_CH1_WIDTH 6
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_RESERVED 31:14
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_XPI_MAP_BITSLIP_WIDTH 14

/* XPI_MAP_CS_OVERRIDE_MASK */
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_OFFSET 16'hee4
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS0 0
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS0_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS1 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS1_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS2 2
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS2_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS3 3
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_PIN_CS3_WIDTH 1
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_RESERVED 31:4
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_FLD_RESERVED_WIDTH 28
`define DDRMC5_MAIN_XPI_MAP_CS_OVERRIDE_MASK_WIDTH 4

/* PAR_ERR_INJ_ECCR */
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_OFFSET 16'hee8
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_SEL0 3:0
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_SEL0_WIDTH 4
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_EN0 4
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_EN0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_DONE0 5
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_DONE0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_PERSISTENT0 6
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_PERSISTENT0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_SEL1 10:7
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_SEL1_WIDTH 4
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_EN1 11
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_EN1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_DONE1 12
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_DONE1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_PERSISTENT1 13
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_PERSISTENT1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAR_ERR_INJ_ECCR_WIDTH 14

/* PAR_ERR_INJ_DBUF */
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_OFFSET 16'heec
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_0 4:0
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_0_WIDTH 5
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_EN0 5
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_EN0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_DONE0 6
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_DONE0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_PERSISTENT0 7
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_PERSISTENT0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_0 12:8
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_0_WIDTH 5
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_EN0 13
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_EN0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_DONE0 14
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_DONE0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_PERSISTENT0 15
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_PERSISTENT0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_1 20:16
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_1_WIDTH 5
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_EN1 21
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_EN1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_DONE1 22
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_DONE1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_PERSISTENT1 23
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_PHY_PERSISTENT1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_1 28:24
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_1_WIDTH 5
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_EN1 29
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_EN1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_DONE1 30
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_DONE1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_PERSISTENT1 31
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_FLD_RAW_PERSISTENT1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_DBUF_WIDTH 32

/* GT_STATUS */
`define DDRMC5_MAIN_GT_STATUS_OFFSET 16'hef0
`define DDRMC5_MAIN_GT_STATUS_FLD_CAPTURE 26:0
`define DDRMC5_MAIN_GT_STATUS_FLD_CAPTURE_WIDTH 27
`define DDRMC5_MAIN_GT_STATUS_FLD_RESERVED 31:27
`define DDRMC5_MAIN_GT_STATUS_FLD_RESERVED_WIDTH 5
`define DDRMC5_MAIN_GT_STATUS_WIDTH 27

/* ALERT_LBDQ_STATUS */
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_OFFSET 16'hef4
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_ALERT 7:0
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_ALERT_WIDTH 8
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_LBDQ 15:8
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_LBDQ_WIDTH 8
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ALERT_LBDQ_STATUS_WIDTH 16

/* ADD_PAR_ERR_INJ */
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_OFFSET 16'hef8
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_PERSISTENT0 0
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_PERSISTENT0_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_SLOT0 2:1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_SLOT0_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_TYPE0 4:3
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_TYPE0_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_EN0 5
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_EN0_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_DONE0 6
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_DONE0_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_CMD0 9:7
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_CMD0_WIDTH 3
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_RANK0 11:10
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_RANK0_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_PERSISTENT1 12
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_PERSISTENT1_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_SLOT1 14:13
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_SLOT1_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_TYPE1 16:15
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_TYPE1_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_EN1 17
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_EN1_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_DONE1 18
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_CMD_DONE1_WIDTH 1
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_CMD1 21:19
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_CMD1_WIDTH 3
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_RANK1 23:22
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_DRAM_RANK1_WIDTH 2
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_RESERVED 31:24
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_ADD_PAR_ERR_INJ_WIDTH 24

/* PAR_ERR_INJ_ILC */
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_OFFSET 16'hefc
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_EN_ILC_0 0
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_EN_ILC_0_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_CTRL_ILC_0 7:1
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_CTRL_ILC_0_WIDTH 7
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_EN_ILC_1 8
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_EN_ILC_1_WIDTH 1
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_CTRL_ILC_1 15:9
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_CTRL_ILC_1_WIDTH 7
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_RESERVED 31:16
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_PAR_ERR_INJ_ILC_WIDTH 16

/* PAR_ERR_LOG_ILC */
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_OFFSET 16'hf00
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_FLD_PAR_ERR_ILC_0 15:0
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_FLD_PAR_ERR_ILC_0_WIDTH 16
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_FLD_PAR_ERR_ILC_1 31:16
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_FLD_PAR_ERR_ILC_1_WIDTH 16
`define DDRMC5_MAIN_PAR_ERR_LOG_ILC_WIDTH 32

/* ILA_CONFIG */
`define DDRMC5_MAIN_ILA_CONFIG_OFFSET 16'hf04
`define DDRMC5_MAIN_ILA_CONFIG_FLD_TRIG_POS 2:0
`define DDRMC5_MAIN_ILA_CONFIG_FLD_TRIG_POS_WIDTH 3
`define DDRMC5_MAIN_ILA_CONFIG_FLD_WINDOW_MASK 10:3
`define DDRMC5_MAIN_ILA_CONFIG_FLD_WINDOW_MASK_WIDTH 8
`define DDRMC5_MAIN_ILA_CONFIG_FLD_TRIG_COND 13:11
`define DDRMC5_MAIN_ILA_CONFIG_FLD_TRIG_COND_WIDTH 3
`define DDRMC5_MAIN_ILA_CONFIG_FLD_HOLD 16:14
`define DDRMC5_MAIN_ILA_CONFIG_FLD_HOLD_WIDTH 3
`define DDRMC5_MAIN_ILA_CONFIG_FLD_RESERVED 31:17
`define DDRMC5_MAIN_ILA_CONFIG_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_ILA_CONFIG_WIDTH 17

/* ILA_STATUS */
`define DDRMC5_MAIN_ILA_STATUS_OFFSET 16'hf08
`define DDRMC5_MAIN_ILA_STATUS_FLD_DONE 0
`define DDRMC5_MAIN_ILA_STATUS_FLD_DONE_WIDTH 1
`define DDRMC5_MAIN_ILA_STATUS_FLD_MATCH 1
`define DDRMC5_MAIN_ILA_STATUS_FLD_MATCH_WIDTH 1
`define DDRMC5_MAIN_ILA_STATUS_FLD_TRIG_SAMPLE 9:2
`define DDRMC5_MAIN_ILA_STATUS_FLD_TRIG_SAMPLE_WIDTH 8
`define DDRMC5_MAIN_ILA_STATUS_FLD_SAMPLE_CNT 17:10
`define DDRMC5_MAIN_ILA_STATUS_FLD_SAMPLE_CNT_WIDTH 8
`define DDRMC5_MAIN_ILA_STATUS_FLD_STATE 20:18
`define DDRMC5_MAIN_ILA_STATUS_FLD_STATE_WIDTH 3
`define DDRMC5_MAIN_ILA_STATUS_FLD_RESERVED 31:21
`define DDRMC5_MAIN_ILA_STATUS_FLD_RESERVED_WIDTH 11
`define DDRMC5_MAIN_ILA_STATUS_WIDTH 21

/* ILA_CAPTURE_DATA */
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_OFFSET 16'hf0c
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_SEL 3:0
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_SEL_WIDTH 4
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_CHANNEL_SEL 4
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_CHANNEL_SEL_WIDTH 1
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_BYTE_SEL 8:5
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_BYTE_SEL_WIDTH 4
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_PHY_NIB_SEL 13:9
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_PHY_NIB_SEL_WIDTH 5
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_OCTAD_SEL 17:14
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_OCTAD_SEL_WIDTH 4
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_DATA_NIB_SEL 21:18
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_DATA_NIB_SEL_WIDTH 4
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_PHASE_SEL 22
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_PHASE_SEL_WIDTH 1
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_CS_SEL 24:23
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_CS_SEL_WIDTH 2
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_RESERVED 31:25
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_FLD_RESERVED_WIDTH 7
`define DDRMC5_MAIN_ILA_CAPTURE_DATA_WIDTH 25

/* ILA_DEBUG_CAL */
`define DDRMC5_MAIN_ILA_DEBUG_CAL_OFFSET 16'hf10
`define DDRMC5_MAIN_ILA_DEBUG_CAL_FLD_SEL 31:0
`define DDRMC5_MAIN_ILA_DEBUG_CAL_FLD_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_DEBUG_CAL_WIDTH 32

/* ILA_CNTRL */
`define DDRMC5_MAIN_ILA_CNTRL_OFFSET 16'hf14
`define DDRMC5_MAIN_ILA_CNTRL_FLD_EN 0
`define DDRMC5_MAIN_ILA_CNTRL_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_ILA_CNTRL_FLD_ARM 1
`define DDRMC5_MAIN_ILA_CNTRL_FLD_ARM_WIDTH 1
`define DDRMC5_MAIN_ILA_CNTRL_FLD_CLK_SEL 2
`define DDRMC5_MAIN_ILA_CNTRL_FLD_CLK_SEL_WIDTH 1
`define DDRMC5_MAIN_ILA_CNTRL_FLD_RESERVED 31:3
`define DDRMC5_MAIN_ILA_CNTRL_FLD_RESERVED_WIDTH 29
`define DDRMC5_MAIN_ILA_CNTRL_WIDTH 3

/* ILA_TRIGGER0 */
`define DDRMC5_MAIN_ILA_TRIGGER0_OFFSET 16'hf18
`define DDRMC5_MAIN_ILA_TRIGGER0_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER0_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER0_WIDTH 32

/* ILA_TRIGGER1 */
`define DDRMC5_MAIN_ILA_TRIGGER1_OFFSET 16'hf1c
`define DDRMC5_MAIN_ILA_TRIGGER1_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER1_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER1_WIDTH 32

/* ILA_TRIGGER2 */
`define DDRMC5_MAIN_ILA_TRIGGER2_OFFSET 16'hf20
`define DDRMC5_MAIN_ILA_TRIGGER2_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER2_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER2_WIDTH 32

/* ILA_TRIGGER3 */
`define DDRMC5_MAIN_ILA_TRIGGER3_OFFSET 16'hf24
`define DDRMC5_MAIN_ILA_TRIGGER3_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER3_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER3_WIDTH 32

/* ILA_TRIGGER4 */
`define DDRMC5_MAIN_ILA_TRIGGER4_OFFSET 16'hf28
`define DDRMC5_MAIN_ILA_TRIGGER4_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER4_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER4_WIDTH 32

/* ILA_TRIGGER5 */
`define DDRMC5_MAIN_ILA_TRIGGER5_OFFSET 16'hf2c
`define DDRMC5_MAIN_ILA_TRIGGER5_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER5_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER5_WIDTH 32

/* ILA_TRIGGER6 */
`define DDRMC5_MAIN_ILA_TRIGGER6_OFFSET 16'hf30
`define DDRMC5_MAIN_ILA_TRIGGER6_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER6_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER6_WIDTH 32

/* ILA_TRIGGER7 */
`define DDRMC5_MAIN_ILA_TRIGGER7_OFFSET 16'hf34
`define DDRMC5_MAIN_ILA_TRIGGER7_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER7_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER7_WIDTH 32

/* ILA_TRIGGER8 */
`define DDRMC5_MAIN_ILA_TRIGGER8_OFFSET 16'hf38
`define DDRMC5_MAIN_ILA_TRIGGER8_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER8_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER8_WIDTH 32

/* ILA_TRIGGER9 */
`define DDRMC5_MAIN_ILA_TRIGGER9_OFFSET 16'hf3c
`define DDRMC5_MAIN_ILA_TRIGGER9_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER9_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER9_WIDTH 32

/* ILA_TRIGGER10 */
`define DDRMC5_MAIN_ILA_TRIGGER10_OFFSET 16'hf40
`define DDRMC5_MAIN_ILA_TRIGGER10_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER10_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER10_WIDTH 32

/* ILA_TRIGGER11 */
`define DDRMC5_MAIN_ILA_TRIGGER11_OFFSET 16'hf44
`define DDRMC5_MAIN_ILA_TRIGGER11_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER11_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER11_WIDTH 32

/* ILA_TRIGGER12 */
`define DDRMC5_MAIN_ILA_TRIGGER12_OFFSET 16'hf48
`define DDRMC5_MAIN_ILA_TRIGGER12_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER12_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER12_WIDTH 32

/* ILA_TRIGGER13 */
`define DDRMC5_MAIN_ILA_TRIGGER13_OFFSET 16'hf4c
`define DDRMC5_MAIN_ILA_TRIGGER13_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER13_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER13_WIDTH 32

/* ILA_TRIGGER14 */
`define DDRMC5_MAIN_ILA_TRIGGER14_OFFSET 16'hf50
`define DDRMC5_MAIN_ILA_TRIGGER14_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER14_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER14_WIDTH 32

/* ILA_TRIGGER15 */
`define DDRMC5_MAIN_ILA_TRIGGER15_OFFSET 16'hf54
`define DDRMC5_MAIN_ILA_TRIGGER15_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER15_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER15_WIDTH 32

/* ILA_TRIGGER16 */
`define DDRMC5_MAIN_ILA_TRIGGER16_OFFSET 16'hf58
`define DDRMC5_MAIN_ILA_TRIGGER16_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER16_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER16_WIDTH 32

/* ILA_TRIGGER17 */
`define DDRMC5_MAIN_ILA_TRIGGER17_OFFSET 16'hf5c
`define DDRMC5_MAIN_ILA_TRIGGER17_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER17_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER17_WIDTH 32

/* ILA_TRIGGER18 */
`define DDRMC5_MAIN_ILA_TRIGGER18_OFFSET 16'hf60
`define DDRMC5_MAIN_ILA_TRIGGER18_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER18_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER18_WIDTH 32

/* ILA_TRIGGER19 */
`define DDRMC5_MAIN_ILA_TRIGGER19_OFFSET 16'hf64
`define DDRMC5_MAIN_ILA_TRIGGER19_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER19_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER19_WIDTH 32

/* ILA_TRIGGER20 */
`define DDRMC5_MAIN_ILA_TRIGGER20_OFFSET 16'hf68
`define DDRMC5_MAIN_ILA_TRIGGER20_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER20_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER20_WIDTH 32

/* ILA_TRIGGER21 */
`define DDRMC5_MAIN_ILA_TRIGGER21_OFFSET 16'hf6c
`define DDRMC5_MAIN_ILA_TRIGGER21_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER21_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER21_WIDTH 32

/* ILA_TRIGGER22 */
`define DDRMC5_MAIN_ILA_TRIGGER22_OFFSET 16'hf70
`define DDRMC5_MAIN_ILA_TRIGGER22_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER22_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER22_WIDTH 32

/* ILA_TRIGGER23 */
`define DDRMC5_MAIN_ILA_TRIGGER23_OFFSET 16'hf74
`define DDRMC5_MAIN_ILA_TRIGGER23_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER23_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER23_WIDTH 32

/* ILA_TRIGGER24 */
`define DDRMC5_MAIN_ILA_TRIGGER24_OFFSET 16'hf78
`define DDRMC5_MAIN_ILA_TRIGGER24_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER24_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER24_WIDTH 32

/* ILA_TRIGGER25 */
`define DDRMC5_MAIN_ILA_TRIGGER25_OFFSET 16'hf7c
`define DDRMC5_MAIN_ILA_TRIGGER25_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER25_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER25_WIDTH 32

/* ILA_TRIGGER26 */
`define DDRMC5_MAIN_ILA_TRIGGER26_OFFSET 16'hf80
`define DDRMC5_MAIN_ILA_TRIGGER26_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER26_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER26_WIDTH 32

/* ILA_TRIGGER27 */
`define DDRMC5_MAIN_ILA_TRIGGER27_OFFSET 16'hf84
`define DDRMC5_MAIN_ILA_TRIGGER27_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER27_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER27_WIDTH 32

/* ILA_TRIGGER28 */
`define DDRMC5_MAIN_ILA_TRIGGER28_OFFSET 16'hf88
`define DDRMC5_MAIN_ILA_TRIGGER28_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER28_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER28_WIDTH 32

/* ILA_TRIGGER29 */
`define DDRMC5_MAIN_ILA_TRIGGER29_OFFSET 16'hf8c
`define DDRMC5_MAIN_ILA_TRIGGER29_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER29_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER29_WIDTH 32

/* ILA_TRIGGER30 */
`define DDRMC5_MAIN_ILA_TRIGGER30_OFFSET 16'hf90
`define DDRMC5_MAIN_ILA_TRIGGER30_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER30_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER30_WIDTH 32

/* ILA_TRIGGER31 */
`define DDRMC5_MAIN_ILA_TRIGGER31_OFFSET 16'hf94
`define DDRMC5_MAIN_ILA_TRIGGER31_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER31_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER31_WIDTH 32

/* ILA_TRIGGER32 */
`define DDRMC5_MAIN_ILA_TRIGGER32_OFFSET 16'hf98
`define DDRMC5_MAIN_ILA_TRIGGER32_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER32_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER32_WIDTH 32

/* ILA_TRIGGER33 */
`define DDRMC5_MAIN_ILA_TRIGGER33_OFFSET 16'hf9c
`define DDRMC5_MAIN_ILA_TRIGGER33_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER33_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER33_WIDTH 32

/* ILA_TRIGGER34 */
`define DDRMC5_MAIN_ILA_TRIGGER34_OFFSET 16'hfa0
`define DDRMC5_MAIN_ILA_TRIGGER34_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER34_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER34_WIDTH 32

/* ILA_TRIGGER35 */
`define DDRMC5_MAIN_ILA_TRIGGER35_OFFSET 16'hfa4
`define DDRMC5_MAIN_ILA_TRIGGER35_FLD_MU 31:0
`define DDRMC5_MAIN_ILA_TRIGGER35_FLD_MU_WIDTH 32
`define DDRMC5_MAIN_ILA_TRIGGER35_WIDTH 32

/* ILA_TRIGGER36 */
`define DDRMC5_MAIN_ILA_TRIGGER36_OFFSET 16'hfa8
`define DDRMC5_MAIN_ILA_TRIGGER36_FLD_MU 8:0
`define DDRMC5_MAIN_ILA_TRIGGER36_FLD_MU_WIDTH 9
`define DDRMC5_MAIN_ILA_TRIGGER36_FLD_RESERVED 31:9
`define DDRMC5_MAIN_ILA_TRIGGER36_FLD_RESERVED_WIDTH 23
`define DDRMC5_MAIN_ILA_TRIGGER36_WIDTH 9

/* ILA_READ_CNTRL */
`define DDRMC5_MAIN_ILA_READ_CNTRL_OFFSET 16'hfac
`define DDRMC5_MAIN_ILA_READ_CNTRL_FLD_ADDR 7:0
`define DDRMC5_MAIN_ILA_READ_CNTRL_FLD_ADDR_WIDTH 8
`define DDRMC5_MAIN_ILA_READ_CNTRL_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ILA_READ_CNTRL_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ILA_READ_CNTRL_WIDTH 8

/* ILA_READ0 */
`define DDRMC5_MAIN_ILA_READ0_OFFSET 16'hfb0
`define DDRMC5_MAIN_ILA_READ0_FLD_DATA 31:0
`define DDRMC5_MAIN_ILA_READ0_FLD_DATA_WIDTH 32
`define DDRMC5_MAIN_ILA_READ0_WIDTH 32

/* ILA_READ1 */
`define DDRMC5_MAIN_ILA_READ1_OFFSET 16'hfb4
`define DDRMC5_MAIN_ILA_READ1_FLD_DATA 31:0
`define DDRMC5_MAIN_ILA_READ1_FLD_DATA_WIDTH 32
`define DDRMC5_MAIN_ILA_READ1_WIDTH 32

/* ILA_READ2 */
`define DDRMC5_MAIN_ILA_READ2_OFFSET 16'hfb8
`define DDRMC5_MAIN_ILA_READ2_FLD_DATA 31:0
`define DDRMC5_MAIN_ILA_READ2_FLD_DATA_WIDTH 32
`define DDRMC5_MAIN_ILA_READ2_WIDTH 32

/* ILA_READ3 */
`define DDRMC5_MAIN_ILA_READ3_OFFSET 16'hfbc
`define DDRMC5_MAIN_ILA_READ3_FLD_DATA 31:0
`define DDRMC5_MAIN_ILA_READ3_FLD_DATA_WIDTH 32
`define DDRMC5_MAIN_ILA_READ3_WIDTH 32

/* ILA_CROSS_TRIG */
`define DDRMC5_MAIN_ILA_CROSS_TRIG_OFFSET 16'hfc0
`define DDRMC5_MAIN_ILA_CROSS_TRIG_FLD_SEL 0
`define DDRMC5_MAIN_ILA_CROSS_TRIG_FLD_SEL_WIDTH 1
`define DDRMC5_MAIN_ILA_CROSS_TRIG_FLD_RESERVED 31:1
`define DDRMC5_MAIN_ILA_CROSS_TRIG_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_ILA_CROSS_TRIG_WIDTH 1

/* DC_PAR_ERR_EN */
`define DDRMC5_MAIN_DC_PAR_ERR_EN_OFFSET 16'hfc4
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_CHK_EN0 0
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_CHK_EN0 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_CHK_EN0 2
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_CHK_EN0 3
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_LOG_EN0 4
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_LOG_EN0 5
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_LOG_EN0 6
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_LOG_EN0 7
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_CHK_EN1 8
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_CHK_EN1 9
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_CHK_EN1 10
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_CHK_EN1 11
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_LOG_EN1 12
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_WBUF2DBUF_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_LOG_EN1 13
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCW_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_LOG_EN1 14
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_DBUF2ECCR_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_LOG_EN1 15
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_ECCR2DBUF_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED 16
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_CHK_EN0 17
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_1 18
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_LOG_EN0 19
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_2 20
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_CHK_EN1 21
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_3 22
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_LOG_EN1 23
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_FARB_ADDR_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_4 31:24
`define DDRMC5_MAIN_DC_PAR_ERR_EN_FLD_RESERVED_4_WIDTH 8
`define DDRMC5_MAIN_DC_PAR_ERR_EN_WIDTH 24

/* DC_ADD_PAR_ERR_LOG0_0 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_0_OFFSET 16'hfc8
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_0_WIDTH 32

/* DC_ADD_PAR_ERR_LOG1_0 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_0_OFFSET 16'hfcc
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_0_WIDTH 32

/* DC_ADD_PAR_ERR_LOG2_0 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_0_OFFSET 16'hfd0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_0_WIDTH 32

/* DC_ADD_PAR_ERR_LOG0_1 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_1_OFFSET 16'hfd4
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG0_1_WIDTH 32

/* DC_ADD_PAR_ERR_LOG1_1 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_1_OFFSET 16'hfd8
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG1_1_WIDTH 32

/* DC_ADD_PAR_ERR_LOG2_1 */
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_1_OFFSET 16'hfdc
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ADD_PAR_ERR_LOG2_1_WIDTH 32

/* DC_DBUF_DATA_PAR_ERR_LOG0_0 */
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_0_OFFSET 16'hfe0
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_0_WIDTH 32

/* DC_DBUF_DATA_PAR_ERR_LOG1_0 */
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_0_OFFSET 16'hfe4
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_0_WIDTH 32

/* DC_DBUF_DATA_PAR_ERR_LOG0_1 */
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_1_OFFSET 16'hfe8
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG0_1_WIDTH 32

/* DC_DBUF_DATA_PAR_ERR_LOG1_1 */
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_1_OFFSET 16'hfec
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_DBUF_DATA_PAR_ERR_LOG1_1_WIDTH 32

/* DC_ECCW_DATA_PAR_ERR_LOG0_0 */
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_0_OFFSET 16'hff0
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_0_WIDTH 32

/* DC_ECCW_DATA_PAR_ERR_LOG0_1 */
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_1_OFFSET 16'hff4
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCW_DATA_PAR_ERR_LOG0_1_WIDTH 32

/* DC_ECCR_DATA_PAR_ERR_LOG0_0 */
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_0_OFFSET 16'hff8
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_0_WIDTH 32

/* DC_ECCR_DATA_PAR_ERR_DATA_LOG0_0 */
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_0_OFFSET 16'hffc
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_0_WIDTH 32

/* DC_ECCR_DATA_PAR_ERR_LOG0_1 */
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_1_OFFSET 16'h1000
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_LOG0_1_WIDTH 32

/* DC_ECCR_DATA_PAR_ERR_DATA_LOG0_1 */
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_1_OFFSET 16'h1004
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_MAIN_DC_ECCR_DATA_PAR_ERR_DATA_LOG0_1_WIDTH 32

/* DC0_PERF_MON */
`define DDRMC5_MAIN_DC0_PERF_MON_OFFSET 16'h1008
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_ENABLE 0
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_ENABLE_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_ACCUM_PERIOD 6:1
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_ACCUM_PERIOD_WIDTH 6
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_NUM_RO 16:7
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_NUM_RO_WIDTH 10
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_NUM_RO_OF 17
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_NUM_RO_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_SNGL 18
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_SNGL_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_DC_ILC_COUNT_SEL 25:19
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_DC_ILC_COUNT_SEL_WIDTH 7
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_RESERVED 31:26
`define DDRMC5_MAIN_DC0_PERF_MON_FLD_RESERVED_WIDTH 6
`define DDRMC5_MAIN_DC0_PERF_MON_WIDTH 26

/* DC0_PERF_MON_ACCU */
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_OFFSET 16'h100c
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_FLD_PERIOD_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_FLD_PERIOD_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_WIDTH 32

/* DC0_PERF_MON_ACCU_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_OFFSET 16'h1010
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_FLD_PERIOD_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_FLD_PERIOD_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_ACCU_HI_WIDTH 16

/* DC0_PERF_MON_0 */
`define DDRMC5_MAIN_DC0_PERF_MON_0_OFFSET 16'h1014
`define DDRMC5_MAIN_DC0_PERF_MON_0_FLD_ACT_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_0_FLD_ACT_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_0_WIDTH 32

/* DC0_PERF_MON_0_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_OFFSET 16'h1018
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_ACT_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_ACT_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_ACT_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_ACT_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_0_HI_WIDTH 17

/* DC0_PERF_MON_1 */
`define DDRMC5_MAIN_DC0_PERF_MON_1_OFFSET 16'h101c
`define DDRMC5_MAIN_DC0_PERF_MON_1_FLD_RD_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_1_FLD_RD_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_1_WIDTH 32

/* DC0_PERF_MON_1_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_OFFSET 16'h1020
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RD_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RD_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RD_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RD_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_1_HI_WIDTH 17

/* DC0_PERF_MON_2 */
`define DDRMC5_MAIN_DC0_PERF_MON_2_OFFSET 16'h1024
`define DDRMC5_MAIN_DC0_PERF_MON_2_FLD_WR_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_2_FLD_WR_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_2_WIDTH 32

/* DC0_PERF_MON_2_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_OFFSET 16'h1028
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_WR_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_WR_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_WR_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_WR_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_2_HI_WIDTH 17

/* DC0_PERF_MON_3 */
`define DDRMC5_MAIN_DC0_PERF_MON_3_OFFSET 16'h102c
`define DDRMC5_MAIN_DC0_PERF_MON_3_FLD_PRE_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_3_FLD_PRE_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_3_WIDTH 32

/* DC0_PERF_MON_3_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_OFFSET 16'h1030
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_PRE_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_PRE_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_PRE_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_PRE_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_3_HI_WIDTH 17

/* DC0_PERF_MON_4 */
`define DDRMC5_MAIN_DC0_PERF_MON_4_OFFSET 16'h1034
`define DDRMC5_MAIN_DC0_PERF_MON_4_FLD_PREA_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_4_FLD_PREA_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_4_WIDTH 32

/* DC0_PERF_MON_4_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_OFFSET 16'h1038
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_PREA_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_PREA_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_PREA_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_PREA_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_4_HI_WIDTH 17

/* DC0_PERF_MON_5 */
`define DDRMC5_MAIN_DC0_PERF_MON_5_OFFSET 16'h103c
`define DDRMC5_MAIN_DC0_PERF_MON_5_FLD_REF_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_5_FLD_REF_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_5_WIDTH 32

/* DC0_PERF_MON_5_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_OFFSET 16'h1040
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_REF_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_REF_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_REF_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_REF_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_5_HI_WIDTH 17

/* DC0_PERF_MON_6 */
`define DDRMC5_MAIN_DC0_PERF_MON_6_OFFSET 16'h1044
`define DDRMC5_MAIN_DC0_PERF_MON_6_FLD_QE_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_6_FLD_QE_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_6_WIDTH 32

/* DC0_PERF_MON_6_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_OFFSET 16'h1048
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_QE_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_QE_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_QE_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_QE_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_6_HI_WIDTH 17

/* DC0_PERF_MON_7 */
`define DDRMC5_MAIN_DC0_PERF_MON_7_OFFSET 16'h104c
`define DDRMC5_MAIN_DC0_PERF_MON_7_FLD_OH_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_7_FLD_OH_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_7_WIDTH 32

/* DC0_PERF_MON_7_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_OFFSET 16'h1050
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_OH_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_OH_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_OH_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_OH_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_7_HI_WIDTH 17

/* DC0_PERF_MON_8 */
`define DDRMC5_MAIN_DC0_PERF_MON_8_OFFSET 16'h1054
`define DDRMC5_MAIN_DC0_PERF_MON_8_FLD_TA_COUNT 31:0
`define DDRMC5_MAIN_DC0_PERF_MON_8_FLD_TA_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC0_PERF_MON_8_WIDTH 32

/* DC0_PERF_MON_8_HI */
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_OFFSET 16'h1058
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_TA_COUNT_HI 15:0
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_TA_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_TA_COUNT_OF 16
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_TA_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC0_PERF_MON_8_HI_WIDTH 17

/* DC1_PERF_MON */
`define DDRMC5_MAIN_DC1_PERF_MON_OFFSET 16'h105c
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_ENABLE 0
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_ENABLE_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_ACCUM_PERIOD 6:1
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_ACCUM_PERIOD_WIDTH 6
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_NUM_RO 16:7
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_NUM_RO_WIDTH 10
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_NUM_RO_OF 17
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_NUM_RO_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_SNGL 18
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_SNGL_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_DC_ILC_COUNT_SEL 25:19
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_DC_ILC_COUNT_SEL_WIDTH 7
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_RESERVED 31:26
`define DDRMC5_MAIN_DC1_PERF_MON_FLD_RESERVED_WIDTH 6
`define DDRMC5_MAIN_DC1_PERF_MON_WIDTH 26

/* DC1_PERF_MON_ACCU */
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_OFFSET 16'h1060
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_FLD_PERIOD_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_FLD_PERIOD_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_WIDTH 32

/* DC1_PERF_MON_ACCU_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_OFFSET 16'h1064
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_FLD_PERIOD_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_FLD_PERIOD_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_ACCU_HI_WIDTH 16

/* DC1_PERF_MON_0 */
`define DDRMC5_MAIN_DC1_PERF_MON_0_OFFSET 16'h1068
`define DDRMC5_MAIN_DC1_PERF_MON_0_FLD_ACT_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_0_FLD_ACT_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_0_WIDTH 32

/* DC1_PERF_MON_0_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_OFFSET 16'h106c
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_ACT_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_ACT_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_ACT_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_ACT_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_0_HI_WIDTH 17

/* DC1_PERF_MON_1 */
`define DDRMC5_MAIN_DC1_PERF_MON_1_OFFSET 16'h1070
`define DDRMC5_MAIN_DC1_PERF_MON_1_FLD_RD_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_1_FLD_RD_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_1_WIDTH 32

/* DC1_PERF_MON_1_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_OFFSET 16'h1074
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RD_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RD_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RD_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RD_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_1_HI_WIDTH 17

/* DC1_PERF_MON_2 */
`define DDRMC5_MAIN_DC1_PERF_MON_2_OFFSET 16'h1078
`define DDRMC5_MAIN_DC1_PERF_MON_2_FLD_WR_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_2_FLD_WR_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_2_WIDTH 32

/* DC1_PERF_MON_2_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_OFFSET 16'h107c
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_WR_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_WR_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_WR_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_WR_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_2_HI_WIDTH 17

/* DC1_PERF_MON_3 */
`define DDRMC5_MAIN_DC1_PERF_MON_3_OFFSET 16'h1080
`define DDRMC5_MAIN_DC1_PERF_MON_3_FLD_PRE_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_3_FLD_PRE_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_3_WIDTH 32

/* DC1_PERF_MON_3_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_OFFSET 16'h1084
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_PRE_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_PRE_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_PRE_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_PRE_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_3_HI_WIDTH 17

/* DC1_PERF_MON_4 */
`define DDRMC5_MAIN_DC1_PERF_MON_4_OFFSET 16'h1088
`define DDRMC5_MAIN_DC1_PERF_MON_4_FLD_PREA_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_4_FLD_PREA_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_4_WIDTH 32

/* DC1_PERF_MON_4_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_OFFSET 16'h108c
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_PREA_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_PREA_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_PREA_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_PREA_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_4_HI_WIDTH 17

/* DC1_PERF_MON_5 */
`define DDRMC5_MAIN_DC1_PERF_MON_5_OFFSET 16'h1090
`define DDRMC5_MAIN_DC1_PERF_MON_5_FLD_REF_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_5_FLD_REF_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_5_WIDTH 32

/* DC1_PERF_MON_5_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_OFFSET 16'h1094
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_REF_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_REF_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_REF_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_REF_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_5_HI_WIDTH 17

/* DC1_PERF_MON_6 */
`define DDRMC5_MAIN_DC1_PERF_MON_6_OFFSET 16'h1098
`define DDRMC5_MAIN_DC1_PERF_MON_6_FLD_QE_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_6_FLD_QE_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_6_WIDTH 32

/* DC1_PERF_MON_6_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_OFFSET 16'h109c
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_QE_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_QE_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_QE_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_QE_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_6_HI_WIDTH 17

/* DC1_PERF_MON_7 */
`define DDRMC5_MAIN_DC1_PERF_MON_7_OFFSET 16'h10a0
`define DDRMC5_MAIN_DC1_PERF_MON_7_FLD_OH_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_7_FLD_OH_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_7_WIDTH 32

/* DC1_PERF_MON_7_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_OFFSET 16'h10a4
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_OH_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_OH_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_OH_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_OH_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_7_HI_WIDTH 17

/* DC1_PERF_MON_8 */
`define DDRMC5_MAIN_DC1_PERF_MON_8_OFFSET 16'h10a8
`define DDRMC5_MAIN_DC1_PERF_MON_8_FLD_TA_COUNT 31:0
`define DDRMC5_MAIN_DC1_PERF_MON_8_FLD_TA_COUNT_WIDTH 32
`define DDRMC5_MAIN_DC1_PERF_MON_8_WIDTH 32

/* DC1_PERF_MON_8_HI */
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_OFFSET 16'h10ac
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_TA_COUNT_HI 15:0
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_TA_COUNT_HI_WIDTH 16
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_TA_COUNT_OF 16
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_TA_COUNT_OF_WIDTH 1
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_RESERVED 31:17
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_DC1_PERF_MON_8_HI_WIDTH 17

/* COMPARE_GT_STATUS_STABLE */
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_OFFSET 16'h10b0
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_FLD_VAL 19:0
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_FLD_VAL_WIDTH 20
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_FLD_RESERVED 31:20
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_COMPARE_GT_STATUS_STABLE_WIDTH 20

/* FIRST_ERR_CAPTURE_ADDR */
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_OFFSET 16'h10b4
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_A 17:0
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_A_WIDTH 18
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_BA 19:18
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_BA_WIDTH 2
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_BG 21:20
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_BG_WIDTH 2
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_RANK 23:22
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_RANK_WIDTH 2
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_CNT 31:24
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_FLD_CNT_WIDTH 8
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_ADDR_WIDTH 32

/* ILA_MUX_D_0_0 */
`define DDRMC5_MAIN_ILA_MUX_D_0_0_OFFSET 16'h10b8
`define DDRMC5_MAIN_ILA_MUX_D_0_0_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_0_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_0_WIDTH 32

/* ILA_MUX_D_0_1 */
`define DDRMC5_MAIN_ILA_MUX_D_0_1_OFFSET 16'h10bc
`define DDRMC5_MAIN_ILA_MUX_D_0_1_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_1_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_1_WIDTH 32

/* ILA_MUX_D_0_2 */
`define DDRMC5_MAIN_ILA_MUX_D_0_2_OFFSET 16'h10c0
`define DDRMC5_MAIN_ILA_MUX_D_0_2_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_2_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_2_WIDTH 32

/* ILA_MUX_D_0_3 */
`define DDRMC5_MAIN_ILA_MUX_D_0_3_OFFSET 16'h10c4
`define DDRMC5_MAIN_ILA_MUX_D_0_3_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_3_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_3_WIDTH 32

/* ILA_MUX_D_0_4 */
`define DDRMC5_MAIN_ILA_MUX_D_0_4_OFFSET 16'h10c8
`define DDRMC5_MAIN_ILA_MUX_D_0_4_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_4_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_4_WIDTH 32

/* ILA_MUX_D_0_5 */
`define DDRMC5_MAIN_ILA_MUX_D_0_5_OFFSET 16'h10cc
`define DDRMC5_MAIN_ILA_MUX_D_0_5_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_5_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_5_WIDTH 32

/* ILA_MUX_D_0_6 */
`define DDRMC5_MAIN_ILA_MUX_D_0_6_OFFSET 16'h10d0
`define DDRMC5_MAIN_ILA_MUX_D_0_6_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_6_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_6_WIDTH 32

/* ILA_MUX_D_0_7 */
`define DDRMC5_MAIN_ILA_MUX_D_0_7_OFFSET 16'h10d4
`define DDRMC5_MAIN_ILA_MUX_D_0_7_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_7_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_7_WIDTH 32

/* ILA_MUX_D_0_8 */
`define DDRMC5_MAIN_ILA_MUX_D_0_8_OFFSET 16'h10d8
`define DDRMC5_MAIN_ILA_MUX_D_0_8_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_8_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_8_WIDTH 32

/* ILA_MUX_D_0_9 */
`define DDRMC5_MAIN_ILA_MUX_D_0_9_OFFSET 16'h10dc
`define DDRMC5_MAIN_ILA_MUX_D_0_9_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_9_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_9_WIDTH 32

/* ILA_MUX_D_0_10 */
`define DDRMC5_MAIN_ILA_MUX_D_0_10_OFFSET 16'h10e0
`define DDRMC5_MAIN_ILA_MUX_D_0_10_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_10_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_10_WIDTH 32

/* ILA_MUX_D_0_11 */
`define DDRMC5_MAIN_ILA_MUX_D_0_11_OFFSET 16'h10e4
`define DDRMC5_MAIN_ILA_MUX_D_0_11_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_11_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_11_WIDTH 32

/* ILA_MUX_D_0_12 */
`define DDRMC5_MAIN_ILA_MUX_D_0_12_OFFSET 16'h10e8
`define DDRMC5_MAIN_ILA_MUX_D_0_12_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_12_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_12_WIDTH 32

/* ILA_MUX_D_0_13 */
`define DDRMC5_MAIN_ILA_MUX_D_0_13_OFFSET 16'h10ec
`define DDRMC5_MAIN_ILA_MUX_D_0_13_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_13_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_13_WIDTH 32

/* ILA_MUX_D_0_14 */
`define DDRMC5_MAIN_ILA_MUX_D_0_14_OFFSET 16'h10f0
`define DDRMC5_MAIN_ILA_MUX_D_0_14_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_14_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_14_WIDTH 32

/* ILA_MUX_D_0_15 */
`define DDRMC5_MAIN_ILA_MUX_D_0_15_OFFSET 16'h10f4
`define DDRMC5_MAIN_ILA_MUX_D_0_15_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_15_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_15_WIDTH 32

/* ILA_MUX_D_0_16 */
`define DDRMC5_MAIN_ILA_MUX_D_0_16_OFFSET 16'h10f8
`define DDRMC5_MAIN_ILA_MUX_D_0_16_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_16_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_16_WIDTH 32

/* ILA_MUX_D_0_17 */
`define DDRMC5_MAIN_ILA_MUX_D_0_17_OFFSET 16'h10fc
`define DDRMC5_MAIN_ILA_MUX_D_0_17_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_0_17_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_0_17_WIDTH 32

/* ILA_MUX_D_1_0 */
`define DDRMC5_MAIN_ILA_MUX_D_1_0_OFFSET 16'h1100
`define DDRMC5_MAIN_ILA_MUX_D_1_0_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_0_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_0_WIDTH 32

/* ILA_MUX_D_1_1 */
`define DDRMC5_MAIN_ILA_MUX_D_1_1_OFFSET 16'h1104
`define DDRMC5_MAIN_ILA_MUX_D_1_1_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_1_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_1_WIDTH 32

/* ILA_MUX_D_1_2 */
`define DDRMC5_MAIN_ILA_MUX_D_1_2_OFFSET 16'h1108
`define DDRMC5_MAIN_ILA_MUX_D_1_2_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_2_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_2_WIDTH 32

/* ILA_MUX_D_1_3 */
`define DDRMC5_MAIN_ILA_MUX_D_1_3_OFFSET 16'h110c
`define DDRMC5_MAIN_ILA_MUX_D_1_3_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_3_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_3_WIDTH 32

/* ILA_MUX_D_1_4 */
`define DDRMC5_MAIN_ILA_MUX_D_1_4_OFFSET 16'h1110
`define DDRMC5_MAIN_ILA_MUX_D_1_4_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_4_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_4_WIDTH 32

/* ILA_MUX_D_1_5 */
`define DDRMC5_MAIN_ILA_MUX_D_1_5_OFFSET 16'h1114
`define DDRMC5_MAIN_ILA_MUX_D_1_5_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_5_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_5_WIDTH 32

/* ILA_MUX_D_1_6 */
`define DDRMC5_MAIN_ILA_MUX_D_1_6_OFFSET 16'h1118
`define DDRMC5_MAIN_ILA_MUX_D_1_6_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_6_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_6_WIDTH 32

/* ILA_MUX_D_1_7 */
`define DDRMC5_MAIN_ILA_MUX_D_1_7_OFFSET 16'h111c
`define DDRMC5_MAIN_ILA_MUX_D_1_7_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_7_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_7_WIDTH 32

/* ILA_MUX_D_1_8 */
`define DDRMC5_MAIN_ILA_MUX_D_1_8_OFFSET 16'h1120
`define DDRMC5_MAIN_ILA_MUX_D_1_8_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_8_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_8_WIDTH 32

/* ILA_MUX_D_1_9 */
`define DDRMC5_MAIN_ILA_MUX_D_1_9_OFFSET 16'h1124
`define DDRMC5_MAIN_ILA_MUX_D_1_9_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_9_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_9_WIDTH 32

/* ILA_MUX_D_1_10 */
`define DDRMC5_MAIN_ILA_MUX_D_1_10_OFFSET 16'h1128
`define DDRMC5_MAIN_ILA_MUX_D_1_10_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_10_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_10_WIDTH 32

/* ILA_MUX_D_1_11 */
`define DDRMC5_MAIN_ILA_MUX_D_1_11_OFFSET 16'h112c
`define DDRMC5_MAIN_ILA_MUX_D_1_11_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_11_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_11_WIDTH 32

/* ILA_MUX_D_1_12 */
`define DDRMC5_MAIN_ILA_MUX_D_1_12_OFFSET 16'h1130
`define DDRMC5_MAIN_ILA_MUX_D_1_12_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_12_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_12_WIDTH 32

/* ILA_MUX_D_1_13 */
`define DDRMC5_MAIN_ILA_MUX_D_1_13_OFFSET 16'h1134
`define DDRMC5_MAIN_ILA_MUX_D_1_13_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_13_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_13_WIDTH 32

/* ILA_MUX_D_1_14 */
`define DDRMC5_MAIN_ILA_MUX_D_1_14_OFFSET 16'h1138
`define DDRMC5_MAIN_ILA_MUX_D_1_14_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_14_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_14_WIDTH 32

/* ILA_MUX_D_1_15 */
`define DDRMC5_MAIN_ILA_MUX_D_1_15_OFFSET 16'h113c
`define DDRMC5_MAIN_ILA_MUX_D_1_15_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_15_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_15_WIDTH 32

/* ILA_MUX_D_1_16 */
`define DDRMC5_MAIN_ILA_MUX_D_1_16_OFFSET 16'h1140
`define DDRMC5_MAIN_ILA_MUX_D_1_16_FLD_DBG_MC_SEL 31:0
`define DDRMC5_MAIN_ILA_MUX_D_1_16_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_MAIN_ILA_MUX_D_1_16_WIDTH 32

/* ILA_MUX_MISC */
`define DDRMC5_MAIN_ILA_MUX_MISC_OFFSET 16'h1144
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_ECCR_DBG_DATA_SEL0 0
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_ECCR_DBG_DATA_SEL0_WIDTH 1
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_ECCR_DBG_DATA_SEL1 1
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_ECCR_DBG_DATA_SEL1_WIDTH 1
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_RESERVED 31:2
`define DDRMC5_MAIN_ILA_MUX_MISC_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_ILA_MUX_MISC_WIDTH 2

/* NOCDBG */
`define DDRMC5_MAIN_NOCDBG_OFFSET 16'h1148
`define DDRMC5_MAIN_NOCDBG_FLD_CLK_SEL 0
`define DDRMC5_MAIN_NOCDBG_FLD_CLK_SEL_WIDTH 1
`define DDRMC5_MAIN_NOCDBG_FLD_CAPTURE_DATA_SEL 3:1
`define DDRMC5_MAIN_NOCDBG_FLD_CAPTURE_DATA_SEL_WIDTH 3
`define DDRMC5_MAIN_NOCDBG_FLD_DATA_DWORD_SEL 5:4
`define DDRMC5_MAIN_NOCDBG_FLD_DATA_DWORD_SEL_WIDTH 2
`define DDRMC5_MAIN_NOCDBG_FLD_RESERVED 31:6
`define DDRMC5_MAIN_NOCDBG_FLD_RESERVED_WIDTH 26
`define DDRMC5_MAIN_NOCDBG_WIDTH 6

/* DDRMC_CLK_CNT */
`define DDRMC5_MAIN_DDRMC_CLK_CNT_OFFSET 16'h114c
`define DDRMC5_MAIN_DDRMC_CLK_CNT_FLD_START_CNT 30:0
`define DDRMC5_MAIN_DDRMC_CLK_CNT_FLD_START_CNT_WIDTH 31
`define DDRMC5_MAIN_DDRMC_CLK_CNT_FLD_START_PULSE 31
`define DDRMC5_MAIN_DDRMC_CLK_CNT_FLD_START_PULSE_WIDTH 1
`define DDRMC5_MAIN_DDRMC_CLK_CNT_WIDTH 32

/* DDRMC_CLK_CNT_STATUS */
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_OFFSET 16'h1150
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_FLD_CURRENT_CNT 30:0
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_FLD_CURRENT_CNT_WIDTH 31
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_FLD_BUSY 31
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_DDRMC_CLK_CNT_STATUS_WIDTH 32

/* PHY_RANK_WRITE_OVERRIDE_DYN */
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_OFFSET 16'h1154
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_ENABLE 1:0
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_ENABLE_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH0_UPDATE_PULSE 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH0_UPDATE_PULSE_WIDTH 1
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH1_UPDATE_PULSE 3
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH1_UPDATE_PULSE_WIDTH 1
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_PAUSE_WRITES 5:4
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_PAUSE_WRITES_WIDTH 2
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH0_RANK_UPDATE 9:6
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH0_RANK_UPDATE_WIDTH 4
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH1_RANK_UPDATE 13:10
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_CH1_RANK_UPDATE_WIDTH 4
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_WRITE_CNT 23:14
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_WRITE_CNT_WIDTH 10
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PHY_RANK_WRITE_OVERRIDE_DYN_WIDTH 24

/* DQI_OSCI_VALUE_LSB_RANK0 */
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_OFFSET 16'h1158
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK0_WIDTH 32

/* DQI_OSCI_VALUE_LSB_RANK1 */
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_OFFSET 16'h115c
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_LSB_RANK1_WIDTH 32

/* DQI_OSCI_VALUE_MSB_RANK0 */
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_OFFSET 16'h1160
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK0_WIDTH 32

/* DQI_OSCI_VALUE_MSB_RANK1 */
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_OFFSET 16'h1164
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQI_OSCI_VALUE_MSB_RANK1_WIDTH 32

/* DQO_OSCI_VALUE_LSB_RANK0 */
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_OFFSET 16'h1168
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK0_WIDTH 32

/* DQO_OSCI_VALUE_LSB_RANK1 */
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_OFFSET 16'h116c
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_LSB_RANK1_WIDTH 32

/* DQO_OSCI_VALUE_MSB_RANK0 */
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_OFFSET 16'h1170
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK0_WIDTH 32

/* DQO_OSCI_VALUE_MSB_RANK1 */
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_OFFSET 16'h1174
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQO_OSCI_VALUE_MSB_RANK1_WIDTH 32

/* DQS_OSCI_VALUE_LSB_0_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_OFFSET 16'h1178
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK0_WIDTH 32

/* DQS_OSCI_VALUE_LSB_1_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_OFFSET 16'h117c
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK0_WIDTH 32

/* DQS_OSCI_VALUE_LSB_2_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_OFFSET 16'h1180
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK0_WIDTH 16

/* DQS_OSCI_VALUE_MSB_0_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_OFFSET 16'h1184
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK0_WIDTH 32

/* DQS_OSCI_VALUE_MSB_1_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_OFFSET 16'h1188
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK0_WIDTH 32

/* DQS_OSCI_VALUE_MSB_2_RANK0 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_OFFSET 16'h118c
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK0_WIDTH 16

/* DQS_OSCI_VALUE_LSB_0_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_OFFSET 16'h1190
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK1_WIDTH 32

/* DQS_OSCI_VALUE_LSB_1_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_OFFSET 16'h1194
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK1_WIDTH 32

/* DQS_OSCI_VALUE_LSB_2_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_OFFSET 16'h1198
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK1_WIDTH 16

/* DQS_OSCI_VALUE_MSB_0_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_OFFSET 16'h119c
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK1_WIDTH 32

/* DQS_OSCI_VALUE_MSB_1_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_OFFSET 16'h11a0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK1_WIDTH 32

/* DQS_OSCI_VALUE_MSB_2_RANK1 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_OFFSET 16'h11a4
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK1_WIDTH 16

/* DQS_OSCI_VALUE_LSB_0_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_OFFSET 16'h11a8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK2_WIDTH 32

/* DQS_OSCI_VALUE_LSB_1_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_OFFSET 16'h11ac
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK2_WIDTH 32

/* DQS_OSCI_VALUE_LSB_2_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_OFFSET 16'h11b0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK2_WIDTH 16

/* DQS_OSCI_VALUE_MSB_0_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_OFFSET 16'h11b4
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK2_WIDTH 32

/* DQS_OSCI_VALUE_MSB_1_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_OFFSET 16'h11b8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK2_WIDTH 32

/* DQS_OSCI_VALUE_MSB_2_RANK2 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_OFFSET 16'h11bc
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK2_WIDTH 16

/* DQS_OSCI_VALUE_LSB_0_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_OFFSET 16'h11c0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_0_RANK3_WIDTH 32

/* DQS_OSCI_VALUE_LSB_1_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_OFFSET 16'h11c4
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_1_RANK3_WIDTH 32

/* DQS_OSCI_VALUE_LSB_2_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_OFFSET 16'h11c8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_LSB_2_RANK3_WIDTH 16

/* DQS_OSCI_VALUE_MSB_0_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_OFFSET 16'h11cc
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_0_RANK3_WIDTH 32

/* DQS_OSCI_VALUE_MSB_1_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_OFFSET 16'h11d0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_1_RANK3_WIDTH 32

/* DQS_OSCI_VALUE_MSB_2_RANK3 */
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_OFFSET 16'h11d4
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DQS_OSCI_VALUE_MSB_2_RANK3_WIDTH 16

/* DRAM_MODE_REG_0 */
`define DDRMC5_MAIN_DRAM_MODE_REG_0_OFFSET 16'h11d8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DRAM_MODE_REG_0_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_0_WIDTH 32

/* DRAM_MODE_REG_1 */
`define DDRMC5_MAIN_DRAM_MODE_REG_1_OFFSET 16'h11dc
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_2 23:16
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_2_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_3 31:24
`define DDRMC5_MAIN_DRAM_MODE_REG_1_FLD_READ_DATA_3_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_1_WIDTH 32

/* DRAM_MODE_REG_2 */
`define DDRMC5_MAIN_DRAM_MODE_REG_2_OFFSET 16'h11e0
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_READ_DATA_0 7:0
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_READ_DATA_0_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_READ_DATA_1 15:8
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_READ_DATA_1_WIDTH 8
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_DRAM_MODE_REG_2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_DRAM_MODE_REG_2_WIDTH 16

/* DRAM_MODE_REG_VALID */
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_OFFSET 16'h11e4
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_CH0 0
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_CH0_WIDTH 1
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_CH1 1
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_CH1_WIDTH 1
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_RESERVED 31:2
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_DRAM_MODE_REG_VALID_WIDTH 2

/* OSCI_STATUS_DDR5_DQS_VALID */
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_OFFSET 16'h11e8
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK0_LSB 0
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK0_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK0_MSB 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK0_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK1_LSB 2
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK1_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK1_MSB 3
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK1_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK2_LSB 4
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK2_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK2_MSB 5
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK2_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK3_LSB 6
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK3_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK3_MSB 7
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RANK3_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RESERVED 31:8
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_OSCI_STATUS_DDR5_DQS_VALID_WIDTH 8

/* OSCI_STATUS_LP5_VALID_CH0 */
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_OFFSET 16'h11ec
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK0_LSB 0
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK0_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK0_MSB 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK0_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK0_LSB 2
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK0_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK0_MSB 3
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK0_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK1_LSB 4
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK1_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK1_MSB 5
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQI_RANK1_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK1_LSB 6
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK1_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK1_MSB 7
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_DQO_RANK1_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_RESERVED 31:8
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH0_WIDTH 8

/* OSCI_STATUS_LP5_VALID_CH1 */
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_OFFSET 16'h11f0
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK0_LSB 0
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK0_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK0_MSB 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK0_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK0_LSB 2
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK0_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK0_MSB 3
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK0_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK1_LSB 4
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK1_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK1_MSB 5
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQI_RANK1_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK1_LSB 6
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK1_LSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK1_MSB 7
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_DQO_RANK1_MSB_WIDTH 1
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_RESERVED 31:8
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_OSCI_STATUS_LP5_VALID_CH1_WIDTH 8

/* MR_READ_ERR_DDR5_OSCI_0 */
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_OFFSET 16'h11f4
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB0 7:0
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB0_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB1 15:8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB1_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB2 23:16
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB2_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB3 31:24
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_FLD_NIB3_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_0_WIDTH 32

/* MR_READ_ERR_DDR5_OSCI_1 */
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_OFFSET 16'h11f8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB4 7:0
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB4_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB5 15:8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB5_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB6 23:16
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB6_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB7 31:24
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_FLD_NIB7_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_1_WIDTH 32

/* MR_READ_ERR_DDR5_OSCI_2 */
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_OFFSET 16'h11fc
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_NIB8 7:0
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_NIB8_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_NIB9 15:8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_NIB9_WIDTH 8
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_OSCI_2_WIDTH 16

/* MR_READ_ERR_DDR5_DRAM_MODE_REG */
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_OFFSET 16'h1200
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_FLD_PER_NIB 9:0
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_FLD_PER_NIB_WIDTH 10
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_FLD_RESERVED 31:10
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_FLD_RESERVED_WIDTH 22
`define DDRMC5_MAIN_MR_READ_ERR_DDR5_DRAM_MODE_REG_WIDTH 10

/* FIRST_ERR_CAPTURE */
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_OFFSET 16'h1204
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_NIBBLE_VALID 17:0
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_NIBBLE_VALID_WIDTH 18
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_BUSY 18
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_FORCE_EN 19
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_FORCE_EN_WIDTH 1
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_RESERVED 31:20
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_FLD_RESERVED_WIDTH 12
`define DDRMC5_MAIN_FIRST_ERR_CAPTURE_WIDTH 20

/* BL16_CAPTURE */
`define DDRMC5_MAIN_BL16_CAPTURE_OFFSET 16'h1208
`define DDRMC5_MAIN_BL16_CAPTURE_FLD_EN 0
`define DDRMC5_MAIN_BL16_CAPTURE_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_BL16_CAPTURE_FLD_RESERVED 31:1
`define DDRMC5_MAIN_BL16_CAPTURE_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_BL16_CAPTURE_WIDTH 1

/* BL16_NIBBLE0 */
`define DDRMC5_MAIN_BL16_NIBBLE0_OFFSET 16'h120c
`define DDRMC5_MAIN_BL16_NIBBLE0_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE0_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE0_WIDTH 32

/* BL16_NIBBLE1 */
`define DDRMC5_MAIN_BL16_NIBBLE1_OFFSET 16'h1210
`define DDRMC5_MAIN_BL16_NIBBLE1_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE1_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE1_WIDTH 32

/* BL16_NIBBLE2 */
`define DDRMC5_MAIN_BL16_NIBBLE2_OFFSET 16'h1214
`define DDRMC5_MAIN_BL16_NIBBLE2_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE2_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE2_WIDTH 32

/* BL16_NIBBLE3 */
`define DDRMC5_MAIN_BL16_NIBBLE3_OFFSET 16'h1218
`define DDRMC5_MAIN_BL16_NIBBLE3_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE3_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE3_WIDTH 32

/* BL16_NIBBLE4 */
`define DDRMC5_MAIN_BL16_NIBBLE4_OFFSET 16'h121c
`define DDRMC5_MAIN_BL16_NIBBLE4_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE4_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE4_WIDTH 32

/* BL16_NIBBLE5 */
`define DDRMC5_MAIN_BL16_NIBBLE5_OFFSET 16'h1220
`define DDRMC5_MAIN_BL16_NIBBLE5_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE5_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE5_WIDTH 32

/* BL16_NIBBLE6 */
`define DDRMC5_MAIN_BL16_NIBBLE6_OFFSET 16'h1224
`define DDRMC5_MAIN_BL16_NIBBLE6_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE6_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE6_WIDTH 32

/* BL16_NIBBLE7 */
`define DDRMC5_MAIN_BL16_NIBBLE7_OFFSET 16'h1228
`define DDRMC5_MAIN_BL16_NIBBLE7_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE7_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE7_WIDTH 32

/* BL16_NIBBLE8 */
`define DDRMC5_MAIN_BL16_NIBBLE8_OFFSET 16'h122c
`define DDRMC5_MAIN_BL16_NIBBLE8_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE8_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE8_WIDTH 32

/* BL16_NIBBLE9 */
`define DDRMC5_MAIN_BL16_NIBBLE9_OFFSET 16'h1230
`define DDRMC5_MAIN_BL16_NIBBLE9_FLD_READ_DATA 31:0
`define DDRMC5_MAIN_BL16_NIBBLE9_FLD_READ_DATA_WIDTH 32
`define DDRMC5_MAIN_BL16_NIBBLE9_WIDTH 32

/* ERR_CNT_NIBBLE0 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_OFFSET 16'h1234
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE0_WIDTH 16

/* ERR_CNT_NIBBLE1 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_OFFSET 16'h1238
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE1_WIDTH 16

/* ERR_CNT_NIBBLE2 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_OFFSET 16'h123c
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE2_WIDTH 16

/* ERR_CNT_NIBBLE3 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_OFFSET 16'h1240
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE3_WIDTH 16

/* ERR_CNT_NIBBLE4 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_OFFSET 16'h1244
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE4_WIDTH 16

/* ERR_CNT_NIBBLE5 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_OFFSET 16'h1248
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE5_WIDTH 16

/* ERR_CNT_NIBBLE6 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_OFFSET 16'h124c
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE6_WIDTH 16

/* ERR_CNT_NIBBLE7 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_OFFSET 16'h1250
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE7_WIDTH 16

/* ERR_CNT_NIBBLE8 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_OFFSET 16'h1254
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE8_WIDTH 16

/* ERR_CNT_NIBBLE9 */
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_OFFSET 16'h1258
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_FLD_VAL 15:0
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ERR_CNT_NIBBLE9_WIDTH 16

/* CPLX_CONFIG */
`define DDRMC5_MAIN_CPLX_CONFIG_OFFSET 16'h125c
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_START 0
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_START_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_WRITE_CAL 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_WRITE_CAL_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_DM_EN 2
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_DM_EN_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_TWOBGBITS_MODE 3
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_TWOBGBITS_MODE_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RANK_EN 7:4
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RANK_EN_WIDTH 4
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_MAX_LOOPS 15:8
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_MAX_LOOPS_WIDTH 8
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_PATTERN_LENGTH 23:16
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_PATTERN_LENGTH_WIDTH 8
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_MAX_BURST_ARRAY_INDEX 28:24
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_MAX_BURST_ARRAY_INDEX_WIDTH 5
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_ISSUE_RESET 29
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_ISSUE_RESET_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RUN_FOREVER 30
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RUN_FOREVER_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RESERVED 31
`define DDRMC5_MAIN_CPLX_CONFIG_FLD_RESERVED_WIDTH 1
`define DDRMC5_MAIN_CPLX_CONFIG_WIDTH 31

/* CPLX_STATUS */
`define DDRMC5_MAIN_CPLX_STATUS_OFFSET 16'h1260
`define DDRMC5_MAIN_CPLX_STATUS_FLD_BUSY 0
`define DDRMC5_MAIN_CPLX_STATUS_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_CPLX_STATUS_FLD_DONE 1
`define DDRMC5_MAIN_CPLX_STATUS_FLD_DONE_WIDTH 1
`define DDRMC5_MAIN_CPLX_STATUS_FLD_RESERVED 31:2
`define DDRMC5_MAIN_CPLX_STATUS_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_CPLX_STATUS_WIDTH 2

/* PRBS_CONFIG */
`define DDRMC5_MAIN_PRBS_CONFIG_OFFSET 16'h1264
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_START 0
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_START_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RD_LOOP 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RD_LOOP_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RUN_FOREVER 2
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RUN_FOREVER_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_ISSUE_RESET 3
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_ISSUE_RESET_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RANK_EN 7:4
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RANK_EN_WIDTH 4
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_REFRESH_EN 8
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_REFRESH_EN_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_DM_EN 9
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_DM_EN_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_TWOBGBITS_MODE 10
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_TWOBGBITS_MODE_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_ONEBABIT_MODE 11
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_ONEBABIT_MODE_WIDTH 1
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_MODE 13:12
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_MODE_WIDTH 2
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_WR_GAP_TIMER_VAL 18:14
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_WR_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RD_GAP_TIMER_VAL 23:19
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RD_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_TWOBGBITSMODE_GAP_TIMER_VAL 28:24
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_TWOBGBITSMODE_GAP_TIMER_VAL_WIDTH 5
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RESERVED 31:29
`define DDRMC5_MAIN_PRBS_CONFIG_FLD_RESERVED_WIDTH 3
`define DDRMC5_MAIN_PRBS_CONFIG_WIDTH 29

/* PRBS_STATUS */
`define DDRMC5_MAIN_PRBS_STATUS_OFFSET 16'h1268
`define DDRMC5_MAIN_PRBS_STATUS_FLD_BUSY 0
`define DDRMC5_MAIN_PRBS_STATUS_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_PRBS_STATUS_FLD_DONE 1
`define DDRMC5_MAIN_PRBS_STATUS_FLD_DONE_WIDTH 1
`define DDRMC5_MAIN_PRBS_STATUS_FLD_RESERVED 31:2
`define DDRMC5_MAIN_PRBS_STATUS_FLD_RESERVED_WIDTH 30
`define DDRMC5_MAIN_PRBS_STATUS_WIDTH 2

/* PRBS_START */
`define DDRMC5_MAIN_PRBS_START_OFFSET 16'h126c
`define DDRMC5_MAIN_PRBS_START_FLD_FLAG 0
`define DDRMC5_MAIN_PRBS_START_FLD_FLAG_WIDTH 1
`define DDRMC5_MAIN_PRBS_START_FLD_RESERVED 31:1
`define DDRMC5_MAIN_PRBS_START_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_PRBS_START_WIDTH 1

/* PAT_DEFAULT_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_OFFSET 16'h1270
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK0_WIDTH 30

/* PAT0_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_OFFSET 16'h1274
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK0_WIDTH 30

/* PAT1_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_OFFSET 16'h1278
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK0_WIDTH 30

/* PAT2_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_OFFSET 16'h127c
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK0_WIDTH 30

/* PAT3_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_OFFSET 16'h1280
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK0_WIDTH 30

/* PAT4_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_OFFSET 16'h1284
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK0_WIDTH 30

/* PAT5_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_OFFSET 16'h1288
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK0_WIDTH 30

/* PAT6_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_OFFSET 16'h128c
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK0_WIDTH 30

/* PAT7_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_OFFSET 16'h1290
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK0_WIDTH 30

/* PAT8_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_OFFSET 16'h1294
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK0_WIDTH 30

/* PAT9_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_OFFSET 16'h1298
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK0_WIDTH 30

/* PAT10_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_OFFSET 16'h129c
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK0_WIDTH 30

/* PAT11_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_OFFSET 16'h12a0
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK0_WIDTH 30

/* PAT12_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_OFFSET 16'h12a4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK0_WIDTH 30

/* PAT13_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_OFFSET 16'h12a8
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK0_WIDTH 30

/* PAT14_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_OFFSET 16'h12ac
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK0_WIDTH 30

/* PAT15_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_OFFSET 16'h12b0
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK0_WIDTH 30

/* PAT16_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_OFFSET 16'h12b4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK0_WIDTH 30

/* PAT17_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_OFFSET 16'h12b8
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK0_WIDTH 30

/* PAT18_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_OFFSET 16'h12bc
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK0_WIDTH 30

/* PAT19_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_OFFSET 16'h12c0
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK0_WIDTH 30

/* PAT20_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_OFFSET 16'h12c4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK0_WIDTH 30

/* PAT21_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_OFFSET 16'h12c8
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK0_WIDTH 30

/* PAT22_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_OFFSET 16'h12cc
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK0_WIDTH 30

/* PAT23_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_OFFSET 16'h12d0
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK0_WIDTH 30

/* PAT24_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_OFFSET 16'h12d4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK0_WIDTH 30

/* PAT25_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_OFFSET 16'h12d8
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK0_WIDTH 30

/* PAT26_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_OFFSET 16'h12dc
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK0_WIDTH 30

/* PAT27_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_OFFSET 16'h12e0
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK0_WIDTH 30

/* PAT28_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_OFFSET 16'h12e4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK0_WIDTH 30

/* PAT29_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_OFFSET 16'h12e8
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK0_WIDTH 30

/* PAT30_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_OFFSET 16'h12ec
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK0_WIDTH 30

/* PAT31_CMD_ADDR_TCK0 */
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_OFFSET 16'h12f0
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA 13:0
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CS 19:16
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CK 26:25
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK0_WIDTH 30

/* PAT_DEFAULT_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_OFFSET 16'h12f4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK1_WIDTH 30

/* PAT0_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_OFFSET 16'h12f8
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK1_WIDTH 30

/* PAT1_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_OFFSET 16'h12fc
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK1_WIDTH 30

/* PAT2_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_OFFSET 16'h1300
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK1_WIDTH 30

/* PAT3_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_OFFSET 16'h1304
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK1_WIDTH 30

/* PAT4_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_OFFSET 16'h1308
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK1_WIDTH 30

/* PAT5_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_OFFSET 16'h130c
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK1_WIDTH 30

/* PAT6_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_OFFSET 16'h1310
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK1_WIDTH 30

/* PAT7_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_OFFSET 16'h1314
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK1_WIDTH 30

/* PAT8_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_OFFSET 16'h1318
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK1_WIDTH 30

/* PAT9_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_OFFSET 16'h131c
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK1_WIDTH 30

/* PAT10_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_OFFSET 16'h1320
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK1_WIDTH 30

/* PAT11_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_OFFSET 16'h1324
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK1_WIDTH 30

/* PAT12_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_OFFSET 16'h1328
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK1_WIDTH 30

/* PAT13_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_OFFSET 16'h132c
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK1_WIDTH 30

/* PAT14_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_OFFSET 16'h1330
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK1_WIDTH 30

/* PAT15_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_OFFSET 16'h1334
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK1_WIDTH 30

/* PAT16_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_OFFSET 16'h1338
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK1_WIDTH 30

/* PAT17_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_OFFSET 16'h133c
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK1_WIDTH 30

/* PAT18_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_OFFSET 16'h1340
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK1_WIDTH 30

/* PAT19_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_OFFSET 16'h1344
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK1_WIDTH 30

/* PAT20_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_OFFSET 16'h1348
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK1_WIDTH 30

/* PAT21_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_OFFSET 16'h134c
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK1_WIDTH 30

/* PAT22_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_OFFSET 16'h1350
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK1_WIDTH 30

/* PAT23_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_OFFSET 16'h1354
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK1_WIDTH 30

/* PAT24_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_OFFSET 16'h1358
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK1_WIDTH 30

/* PAT25_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_OFFSET 16'h135c
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK1_WIDTH 30

/* PAT26_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_OFFSET 16'h1360
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK1_WIDTH 30

/* PAT27_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_OFFSET 16'h1364
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK1_WIDTH 30

/* PAT28_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_OFFSET 16'h1368
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK1_WIDTH 30

/* PAT29_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_OFFSET 16'h136c
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK1_WIDTH 30

/* PAT30_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_OFFSET 16'h1370
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK1_WIDTH 30

/* PAT31_CMD_ADDR_TCK1 */
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_OFFSET 16'h1374
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA 13:0
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CS 19:16
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CK 26:25
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK1_WIDTH 30

/* PAT_DEFAULT_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_OFFSET 16'h1378
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK2_WIDTH 30

/* PAT0_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_OFFSET 16'h137c
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK2_WIDTH 30

/* PAT1_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_OFFSET 16'h1380
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK2_WIDTH 30

/* PAT2_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_OFFSET 16'h1384
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK2_WIDTH 30

/* PAT3_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_OFFSET 16'h1388
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK2_WIDTH 30

/* PAT4_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_OFFSET 16'h138c
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK2_WIDTH 30

/* PAT5_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_OFFSET 16'h1390
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK2_WIDTH 30

/* PAT6_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_OFFSET 16'h1394
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK2_WIDTH 30

/* PAT7_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_OFFSET 16'h1398
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK2_WIDTH 30

/* PAT8_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_OFFSET 16'h139c
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK2_WIDTH 30

/* PAT9_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_OFFSET 16'h13a0
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK2_WIDTH 30

/* PAT10_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_OFFSET 16'h13a4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK2_WIDTH 30

/* PAT11_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_OFFSET 16'h13a8
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK2_WIDTH 30

/* PAT12_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_OFFSET 16'h13ac
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK2_WIDTH 30

/* PAT13_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_OFFSET 16'h13b0
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK2_WIDTH 30

/* PAT14_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_OFFSET 16'h13b4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK2_WIDTH 30

/* PAT15_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_OFFSET 16'h13b8
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK2_WIDTH 30

/* PAT16_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_OFFSET 16'h13bc
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK2_WIDTH 30

/* PAT17_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_OFFSET 16'h13c0
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK2_WIDTH 30

/* PAT18_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_OFFSET 16'h13c4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK2_WIDTH 30

/* PAT19_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_OFFSET 16'h13c8
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK2_WIDTH 30

/* PAT20_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_OFFSET 16'h13cc
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK2_WIDTH 30

/* PAT21_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_OFFSET 16'h13d0
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK2_WIDTH 30

/* PAT22_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_OFFSET 16'h13d4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK2_WIDTH 30

/* PAT23_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_OFFSET 16'h13d8
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK2_WIDTH 30

/* PAT24_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_OFFSET 16'h13dc
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK2_WIDTH 30

/* PAT25_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_OFFSET 16'h13e0
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK2_WIDTH 30

/* PAT26_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_OFFSET 16'h13e4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK2_WIDTH 30

/* PAT27_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_OFFSET 16'h13e8
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK2_WIDTH 30

/* PAT28_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_OFFSET 16'h13ec
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK2_WIDTH 30

/* PAT29_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_OFFSET 16'h13f0
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK2_WIDTH 30

/* PAT30_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_OFFSET 16'h13f4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK2_WIDTH 30

/* PAT31_CMD_ADDR_TCK2 */
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_OFFSET 16'h13f8
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA 13:0
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CS 19:16
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CK 26:25
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK2_WIDTH 30

/* PAT_DEFAULT_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_OFFSET 16'h13fc
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT_DEFAULT_CMD_ADDR_TCK3_WIDTH 30

/* PAT0_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_OFFSET 16'h1400
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT0_CMD_ADDR_TCK3_WIDTH 30

/* PAT1_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_OFFSET 16'h1404
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT1_CMD_ADDR_TCK3_WIDTH 30

/* PAT2_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_OFFSET 16'h1408
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT2_CMD_ADDR_TCK3_WIDTH 30

/* PAT3_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_OFFSET 16'h140c
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT3_CMD_ADDR_TCK3_WIDTH 30

/* PAT4_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_OFFSET 16'h1410
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT4_CMD_ADDR_TCK3_WIDTH 30

/* PAT5_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_OFFSET 16'h1414
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT5_CMD_ADDR_TCK3_WIDTH 30

/* PAT6_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_OFFSET 16'h1418
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT6_CMD_ADDR_TCK3_WIDTH 30

/* PAT7_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_OFFSET 16'h141c
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT7_CMD_ADDR_TCK3_WIDTH 30

/* PAT8_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_OFFSET 16'h1420
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT8_CMD_ADDR_TCK3_WIDTH 30

/* PAT9_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_OFFSET 16'h1424
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT9_CMD_ADDR_TCK3_WIDTH 30

/* PAT10_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_OFFSET 16'h1428
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT10_CMD_ADDR_TCK3_WIDTH 30

/* PAT11_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_OFFSET 16'h142c
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT11_CMD_ADDR_TCK3_WIDTH 30

/* PAT12_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_OFFSET 16'h1430
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT12_CMD_ADDR_TCK3_WIDTH 30

/* PAT13_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_OFFSET 16'h1434
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT13_CMD_ADDR_TCK3_WIDTH 30

/* PAT14_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_OFFSET 16'h1438
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT14_CMD_ADDR_TCK3_WIDTH 30

/* PAT15_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_OFFSET 16'h143c
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT15_CMD_ADDR_TCK3_WIDTH 30

/* PAT16_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_OFFSET 16'h1440
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT16_CMD_ADDR_TCK3_WIDTH 30

/* PAT17_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_OFFSET 16'h1444
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT17_CMD_ADDR_TCK3_WIDTH 30

/* PAT18_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_OFFSET 16'h1448
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT18_CMD_ADDR_TCK3_WIDTH 30

/* PAT19_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_OFFSET 16'h144c
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT19_CMD_ADDR_TCK3_WIDTH 30

/* PAT20_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_OFFSET 16'h1450
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT20_CMD_ADDR_TCK3_WIDTH 30

/* PAT21_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_OFFSET 16'h1454
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT21_CMD_ADDR_TCK3_WIDTH 30

/* PAT22_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_OFFSET 16'h1458
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT22_CMD_ADDR_TCK3_WIDTH 30

/* PAT23_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_OFFSET 16'h145c
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT23_CMD_ADDR_TCK3_WIDTH 30

/* PAT24_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_OFFSET 16'h1460
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT24_CMD_ADDR_TCK3_WIDTH 30

/* PAT25_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_OFFSET 16'h1464
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT25_CMD_ADDR_TCK3_WIDTH 30

/* PAT26_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_OFFSET 16'h1468
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT26_CMD_ADDR_TCK3_WIDTH 30

/* PAT27_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_OFFSET 16'h146c
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT27_CMD_ADDR_TCK3_WIDTH 30

/* PAT28_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_OFFSET 16'h1470
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT28_CMD_ADDR_TCK3_WIDTH 30

/* PAT29_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_OFFSET 16'h1474
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT29_CMD_ADDR_TCK3_WIDTH 30

/* PAT30_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_OFFSET 16'h1478
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT30_CMD_ADDR_TCK3_WIDTH 30

/* PAT31_CMD_ADDR_TCK3 */
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_OFFSET 16'h147c
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA 13:0
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_WIDTH 14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_PAR 15:14
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_PAR_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CS 19:16
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS 23:20
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_INC_DEC_BIT_POS_WIDTH 4
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_RESET_N 24
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_RESET_N_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CK 26:25
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CK_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE 27
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_TYPE_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC 28
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_SRC_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN 29
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_CA_UPDATE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_RESERVED 31:30
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_FLD_RESERVED_WIDTH 2
`define DDRMC5_MAIN_PAT31_CMD_ADDR_TCK3_WIDTH 30

/* PAT_DEFAULT_CAS */
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_OFFSET 16'h1480
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT_DEFAULT_CAS_WIDTH 13

/* PAT0_CAS */
`define DDRMC5_MAIN_PAT0_CAS_OFFSET 16'h1484
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT0_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT0_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT0_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT0_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT0_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT0_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT0_CAS_WIDTH 13

/* PAT1_CAS */
`define DDRMC5_MAIN_PAT1_CAS_OFFSET 16'h1488
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT1_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT1_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT1_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT1_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT1_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT1_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT1_CAS_WIDTH 13

/* PAT2_CAS */
`define DDRMC5_MAIN_PAT2_CAS_OFFSET 16'h148c
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT2_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT2_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT2_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT2_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT2_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT2_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT2_CAS_WIDTH 13

/* PAT3_CAS */
`define DDRMC5_MAIN_PAT3_CAS_OFFSET 16'h1490
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT3_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT3_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT3_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT3_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT3_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT3_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT3_CAS_WIDTH 13

/* PAT4_CAS */
`define DDRMC5_MAIN_PAT4_CAS_OFFSET 16'h1494
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT4_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT4_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT4_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT4_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT4_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT4_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT4_CAS_WIDTH 13

/* PAT5_CAS */
`define DDRMC5_MAIN_PAT5_CAS_OFFSET 16'h1498
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT5_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT5_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT5_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT5_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT5_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT5_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT5_CAS_WIDTH 13

/* PAT6_CAS */
`define DDRMC5_MAIN_PAT6_CAS_OFFSET 16'h149c
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT6_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT6_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT6_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT6_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT6_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT6_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT6_CAS_WIDTH 13

/* PAT7_CAS */
`define DDRMC5_MAIN_PAT7_CAS_OFFSET 16'h14a0
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT7_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT7_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT7_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT7_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT7_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT7_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT7_CAS_WIDTH 13

/* PAT8_CAS */
`define DDRMC5_MAIN_PAT8_CAS_OFFSET 16'h14a4
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT8_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT8_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT8_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT8_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT8_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT8_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT8_CAS_WIDTH 13

/* PAT9_CAS */
`define DDRMC5_MAIN_PAT9_CAS_OFFSET 16'h14a8
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT9_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT9_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT9_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT9_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT9_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT9_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT9_CAS_WIDTH 13

/* PAT10_CAS */
`define DDRMC5_MAIN_PAT10_CAS_OFFSET 16'h14ac
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT10_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT10_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT10_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT10_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT10_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT10_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT10_CAS_WIDTH 13

/* PAT11_CAS */
`define DDRMC5_MAIN_PAT11_CAS_OFFSET 16'h14b0
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT11_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT11_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT11_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT11_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT11_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT11_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT11_CAS_WIDTH 13

/* PAT12_CAS */
`define DDRMC5_MAIN_PAT12_CAS_OFFSET 16'h14b4
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT12_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT12_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT12_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT12_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT12_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT12_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT12_CAS_WIDTH 13

/* PAT13_CAS */
`define DDRMC5_MAIN_PAT13_CAS_OFFSET 16'h14b8
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT13_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT13_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT13_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT13_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT13_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT13_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT13_CAS_WIDTH 13

/* PAT14_CAS */
`define DDRMC5_MAIN_PAT14_CAS_OFFSET 16'h14bc
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT14_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT14_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT14_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT14_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT14_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT14_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT14_CAS_WIDTH 13

/* PAT15_CAS */
`define DDRMC5_MAIN_PAT15_CAS_OFFSET 16'h14c0
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT15_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT15_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT15_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT15_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT15_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT15_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT15_CAS_WIDTH 13

/* PAT16_CAS */
`define DDRMC5_MAIN_PAT16_CAS_OFFSET 16'h14c4
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT16_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT16_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT16_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT16_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT16_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT16_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT16_CAS_WIDTH 13

/* PAT17_CAS */
`define DDRMC5_MAIN_PAT17_CAS_OFFSET 16'h14c8
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT17_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT17_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT17_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT17_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT17_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT17_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT17_CAS_WIDTH 13

/* PAT18_CAS */
`define DDRMC5_MAIN_PAT18_CAS_OFFSET 16'h14cc
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT18_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT18_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT18_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT18_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT18_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT18_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT18_CAS_WIDTH 13

/* PAT19_CAS */
`define DDRMC5_MAIN_PAT19_CAS_OFFSET 16'h14d0
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT19_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT19_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT19_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT19_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT19_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT19_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT19_CAS_WIDTH 13

/* PAT20_CAS */
`define DDRMC5_MAIN_PAT20_CAS_OFFSET 16'h14d4
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT20_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT20_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT20_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT20_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT20_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT20_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT20_CAS_WIDTH 13

/* PAT21_CAS */
`define DDRMC5_MAIN_PAT21_CAS_OFFSET 16'h14d8
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT21_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT21_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT21_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT21_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT21_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT21_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT21_CAS_WIDTH 13

/* PAT22_CAS */
`define DDRMC5_MAIN_PAT22_CAS_OFFSET 16'h14dc
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT22_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT22_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT22_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT22_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT22_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT22_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT22_CAS_WIDTH 13

/* PAT23_CAS */
`define DDRMC5_MAIN_PAT23_CAS_OFFSET 16'h14e0
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT23_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT23_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT23_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT23_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT23_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT23_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT23_CAS_WIDTH 13

/* PAT24_CAS */
`define DDRMC5_MAIN_PAT24_CAS_OFFSET 16'h14e4
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT24_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT24_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT24_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT24_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT24_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT24_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT24_CAS_WIDTH 13

/* PAT25_CAS */
`define DDRMC5_MAIN_PAT25_CAS_OFFSET 16'h14e8
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT25_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT25_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT25_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT25_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT25_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT25_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT25_CAS_WIDTH 13

/* PAT26_CAS */
`define DDRMC5_MAIN_PAT26_CAS_OFFSET 16'h14ec
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT26_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT26_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT26_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT26_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT26_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT26_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT26_CAS_WIDTH 13

/* PAT27_CAS */
`define DDRMC5_MAIN_PAT27_CAS_OFFSET 16'h14f0
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT27_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT27_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT27_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT27_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT27_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT27_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT27_CAS_WIDTH 13

/* PAT28_CAS */
`define DDRMC5_MAIN_PAT28_CAS_OFFSET 16'h14f4
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT28_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT28_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT28_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT28_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT28_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT28_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT28_CAS_WIDTH 13

/* PAT29_CAS */
`define DDRMC5_MAIN_PAT29_CAS_OFFSET 16'h14f8
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT29_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT29_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT29_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT29_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT29_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT29_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT29_CAS_WIDTH 13

/* PAT30_CAS */
`define DDRMC5_MAIN_PAT30_CAS_OFFSET 16'h14fc
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT30_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT30_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT30_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT30_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT30_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT30_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT30_CAS_WIDTH 13

/* PAT31_CAS */
`define DDRMC5_MAIN_PAT31_CAS_OFFSET 16'h1500
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK0 0
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK0 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK1 2
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK1 3
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK2 4
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK2 5
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK3 6
`define DDRMC5_MAIN_PAT31_CAS_FLD_EN_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK3 7
`define DDRMC5_MAIN_PAT31_CAS_FLD_RD_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK0 8
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK1 9
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK2 10
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK3 11
`define DDRMC5_MAIN_PAT31_CAS_FLD_WS_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_CA_DRIVE_DISABLE 12
`define DDRMC5_MAIN_PAT31_CAS_FLD_CA_DRIVE_DISABLE_WIDTH 1
`define DDRMC5_MAIN_PAT31_CAS_FLD_RESERVED 31:13
`define DDRMC5_MAIN_PAT31_CAS_FLD_RESERVED_WIDTH 19
`define DDRMC5_MAIN_PAT31_CAS_WIDTH 13

/* PAT_DEFAULT_DQ */
`define DDRMC5_MAIN_PAT_DEFAULT_DQ_OFFSET 16'h1504
`define DDRMC5_MAIN_PAT_DEFAULT_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT_DEFAULT_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT_DEFAULT_DQ_WIDTH 32

/* PAT0_DQ */
`define DDRMC5_MAIN_PAT0_DQ_OFFSET 16'h1508
`define DDRMC5_MAIN_PAT0_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT0_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT0_DQ_WIDTH 32

/* PAT1_DQ */
`define DDRMC5_MAIN_PAT1_DQ_OFFSET 16'h150c
`define DDRMC5_MAIN_PAT1_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT1_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT1_DQ_WIDTH 32

/* PAT2_DQ */
`define DDRMC5_MAIN_PAT2_DQ_OFFSET 16'h1510
`define DDRMC5_MAIN_PAT2_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT2_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT2_DQ_WIDTH 32

/* PAT3_DQ */
`define DDRMC5_MAIN_PAT3_DQ_OFFSET 16'h1514
`define DDRMC5_MAIN_PAT3_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT3_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT3_DQ_WIDTH 32

/* PAT4_DQ */
`define DDRMC5_MAIN_PAT4_DQ_OFFSET 16'h1518
`define DDRMC5_MAIN_PAT4_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT4_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT4_DQ_WIDTH 32

/* PAT5_DQ */
`define DDRMC5_MAIN_PAT5_DQ_OFFSET 16'h151c
`define DDRMC5_MAIN_PAT5_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT5_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT5_DQ_WIDTH 32

/* PAT6_DQ */
`define DDRMC5_MAIN_PAT6_DQ_OFFSET 16'h1520
`define DDRMC5_MAIN_PAT6_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT6_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT6_DQ_WIDTH 32

/* PAT7_DQ */
`define DDRMC5_MAIN_PAT7_DQ_OFFSET 16'h1524
`define DDRMC5_MAIN_PAT7_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT7_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT7_DQ_WIDTH 32

/* PAT8_DQ */
`define DDRMC5_MAIN_PAT8_DQ_OFFSET 16'h1528
`define DDRMC5_MAIN_PAT8_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT8_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT8_DQ_WIDTH 32

/* PAT9_DQ */
`define DDRMC5_MAIN_PAT9_DQ_OFFSET 16'h152c
`define DDRMC5_MAIN_PAT9_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT9_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT9_DQ_WIDTH 32

/* PAT10_DQ */
`define DDRMC5_MAIN_PAT10_DQ_OFFSET 16'h1530
`define DDRMC5_MAIN_PAT10_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT10_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT10_DQ_WIDTH 32

/* PAT11_DQ */
`define DDRMC5_MAIN_PAT11_DQ_OFFSET 16'h1534
`define DDRMC5_MAIN_PAT11_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT11_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT11_DQ_WIDTH 32

/* PAT12_DQ */
`define DDRMC5_MAIN_PAT12_DQ_OFFSET 16'h1538
`define DDRMC5_MAIN_PAT12_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT12_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT12_DQ_WIDTH 32

/* PAT13_DQ */
`define DDRMC5_MAIN_PAT13_DQ_OFFSET 16'h153c
`define DDRMC5_MAIN_PAT13_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT13_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT13_DQ_WIDTH 32

/* PAT14_DQ */
`define DDRMC5_MAIN_PAT14_DQ_OFFSET 16'h1540
`define DDRMC5_MAIN_PAT14_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT14_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT14_DQ_WIDTH 32

/* PAT15_DQ */
`define DDRMC5_MAIN_PAT15_DQ_OFFSET 16'h1544
`define DDRMC5_MAIN_PAT15_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT15_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT15_DQ_WIDTH 32

/* PAT16_DQ */
`define DDRMC5_MAIN_PAT16_DQ_OFFSET 16'h1548
`define DDRMC5_MAIN_PAT16_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT16_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT16_DQ_WIDTH 32

/* PAT17_DQ */
`define DDRMC5_MAIN_PAT17_DQ_OFFSET 16'h154c
`define DDRMC5_MAIN_PAT17_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT17_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT17_DQ_WIDTH 32

/* PAT18_DQ */
`define DDRMC5_MAIN_PAT18_DQ_OFFSET 16'h1550
`define DDRMC5_MAIN_PAT18_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT18_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT18_DQ_WIDTH 32

/* PAT19_DQ */
`define DDRMC5_MAIN_PAT19_DQ_OFFSET 16'h1554
`define DDRMC5_MAIN_PAT19_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT19_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT19_DQ_WIDTH 32

/* PAT20_DQ */
`define DDRMC5_MAIN_PAT20_DQ_OFFSET 16'h1558
`define DDRMC5_MAIN_PAT20_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT20_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT20_DQ_WIDTH 32

/* PAT21_DQ */
`define DDRMC5_MAIN_PAT21_DQ_OFFSET 16'h155c
`define DDRMC5_MAIN_PAT21_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT21_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT21_DQ_WIDTH 32

/* PAT22_DQ */
`define DDRMC5_MAIN_PAT22_DQ_OFFSET 16'h1560
`define DDRMC5_MAIN_PAT22_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT22_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT22_DQ_WIDTH 32

/* PAT23_DQ */
`define DDRMC5_MAIN_PAT23_DQ_OFFSET 16'h1564
`define DDRMC5_MAIN_PAT23_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT23_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT23_DQ_WIDTH 32

/* PAT24_DQ */
`define DDRMC5_MAIN_PAT24_DQ_OFFSET 16'h1568
`define DDRMC5_MAIN_PAT24_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT24_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT24_DQ_WIDTH 32

/* PAT25_DQ */
`define DDRMC5_MAIN_PAT25_DQ_OFFSET 16'h156c
`define DDRMC5_MAIN_PAT25_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT25_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT25_DQ_WIDTH 32

/* PAT26_DQ */
`define DDRMC5_MAIN_PAT26_DQ_OFFSET 16'h1570
`define DDRMC5_MAIN_PAT26_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT26_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT26_DQ_WIDTH 32

/* PAT27_DQ */
`define DDRMC5_MAIN_PAT27_DQ_OFFSET 16'h1574
`define DDRMC5_MAIN_PAT27_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT27_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT27_DQ_WIDTH 32

/* PAT28_DQ */
`define DDRMC5_MAIN_PAT28_DQ_OFFSET 16'h1578
`define DDRMC5_MAIN_PAT28_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT28_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT28_DQ_WIDTH 32

/* PAT29_DQ */
`define DDRMC5_MAIN_PAT29_DQ_OFFSET 16'h157c
`define DDRMC5_MAIN_PAT29_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT29_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT29_DQ_WIDTH 32

/* PAT30_DQ */
`define DDRMC5_MAIN_PAT30_DQ_OFFSET 16'h1580
`define DDRMC5_MAIN_PAT30_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT30_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT30_DQ_WIDTH 32

/* PAT31_DQ */
`define DDRMC5_MAIN_PAT31_DQ_OFFSET 16'h1584
`define DDRMC5_MAIN_PAT31_DQ_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT31_DQ_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT31_DQ_WIDTH 32

/* PAT_DEFAULT_DMDBI_DQS */
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_OFFSET 16'h1588
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT_DEFAULT_DMDBI_DQS_WIDTH 24

/* PAT0_DMDBI_DQS */
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_OFFSET 16'h158c
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT0_DMDBI_DQS_WIDTH 24

/* PAT1_DMDBI_DQS */
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_OFFSET 16'h1590
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT1_DMDBI_DQS_WIDTH 24

/* PAT2_DMDBI_DQS */
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_OFFSET 16'h1594
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT2_DMDBI_DQS_WIDTH 24

/* PAT3_DMDBI_DQS */
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_OFFSET 16'h1598
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT3_DMDBI_DQS_WIDTH 24

/* PAT4_DMDBI_DQS */
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_OFFSET 16'h159c
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT4_DMDBI_DQS_WIDTH 24

/* PAT5_DMDBI_DQS */
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_OFFSET 16'h15a0
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT5_DMDBI_DQS_WIDTH 24

/* PAT6_DMDBI_DQS */
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_OFFSET 16'h15a4
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT6_DMDBI_DQS_WIDTH 24

/* PAT7_DMDBI_DQS */
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_OFFSET 16'h15a8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT7_DMDBI_DQS_WIDTH 24

/* PAT8_DMDBI_DQS */
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_OFFSET 16'h15ac
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT8_DMDBI_DQS_WIDTH 24

/* PAT9_DMDBI_DQS */
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_OFFSET 16'h15b0
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT9_DMDBI_DQS_WIDTH 24

/* PAT10_DMDBI_DQS */
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_OFFSET 16'h15b4
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT10_DMDBI_DQS_WIDTH 24

/* PAT11_DMDBI_DQS */
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_OFFSET 16'h15b8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT11_DMDBI_DQS_WIDTH 24

/* PAT12_DMDBI_DQS */
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_OFFSET 16'h15bc
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT12_DMDBI_DQS_WIDTH 24

/* PAT13_DMDBI_DQS */
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_OFFSET 16'h15c0
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT13_DMDBI_DQS_WIDTH 24

/* PAT14_DMDBI_DQS */
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_OFFSET 16'h15c4
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT14_DMDBI_DQS_WIDTH 24

/* PAT15_DMDBI_DQS */
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_OFFSET 16'h15c8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT15_DMDBI_DQS_WIDTH 24

/* PAT16_DMDBI_DQS */
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_OFFSET 16'h15cc
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT16_DMDBI_DQS_WIDTH 24

/* PAT17_DMDBI_DQS */
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_OFFSET 16'h15d0
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT17_DMDBI_DQS_WIDTH 24

/* PAT18_DMDBI_DQS */
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_OFFSET 16'h15d4
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT18_DMDBI_DQS_WIDTH 24

/* PAT19_DMDBI_DQS */
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_OFFSET 16'h15d8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT19_DMDBI_DQS_WIDTH 24

/* PAT20_DMDBI_DQS */
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_OFFSET 16'h15dc
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT20_DMDBI_DQS_WIDTH 24

/* PAT21_DMDBI_DQS */
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_OFFSET 16'h15e0
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT21_DMDBI_DQS_WIDTH 24

/* PAT22_DMDBI_DQS */
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_OFFSET 16'h15e4
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT22_DMDBI_DQS_WIDTH 24

/* PAT23_DMDBI_DQS */
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_OFFSET 16'h15e8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT23_DMDBI_DQS_WIDTH 24

/* PAT24_DMDBI_DQS */
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_OFFSET 16'h15ec
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT24_DMDBI_DQS_WIDTH 24

/* PAT25_DMDBI_DQS */
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_OFFSET 16'h15f0
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT25_DMDBI_DQS_WIDTH 24

/* PAT26_DMDBI_DQS */
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_OFFSET 16'h15f4
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT26_DMDBI_DQS_WIDTH 24

/* PAT27_DMDBI_DQS */
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_OFFSET 16'h15f8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT27_DMDBI_DQS_WIDTH 24

/* PAT28_DMDBI_DQS */
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_OFFSET 16'h15fc
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT28_DMDBI_DQS_WIDTH 24

/* PAT29_DMDBI_DQS */
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_OFFSET 16'h1600
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT29_DMDBI_DQS_WIDTH 24

/* PAT30_DMDBI_DQS */
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_OFFSET 16'h1604
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT30_DMDBI_DQS_WIDTH 24

/* PAT31_DMDBI_DQS */
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_OFFSET 16'h1608
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_DMDBI 7:0
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_DMDBI_WIDTH 8
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_DQS 15:8
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_DQS_WIDTH 8
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_EDGE_CMPR_MASK 23:16
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_EDGE_CMPR_MASK_WIDTH 8
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_RESERVED 31:24
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_FLD_RESERVED_WIDTH 8
`define DDRMC5_MAIN_PAT31_DMDBI_DQS_WIDTH 24

/* DEFAULT_PAT_EXE_CFG_INNER */
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_OFFSET 16'h160c
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_INNER_WIDTH 32

/* PAT0_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_OFFSET 16'h1610
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT0_EXE_CFG_INNER_WIDTH 32

/* PAT1_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_OFFSET 16'h1614
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT1_EXE_CFG_INNER_WIDTH 32

/* PAT2_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_OFFSET 16'h1618
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT2_EXE_CFG_INNER_WIDTH 32

/* PAT3_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_OFFSET 16'h161c
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT3_EXE_CFG_INNER_WIDTH 32

/* PAT4_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_OFFSET 16'h1620
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT4_EXE_CFG_INNER_WIDTH 32

/* PAT5_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_OFFSET 16'h1624
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT5_EXE_CFG_INNER_WIDTH 32

/* PAT6_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_OFFSET 16'h1628
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT6_EXE_CFG_INNER_WIDTH 32

/* PAT7_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_OFFSET 16'h162c
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT7_EXE_CFG_INNER_WIDTH 32

/* PAT8_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_OFFSET 16'h1630
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT8_EXE_CFG_INNER_WIDTH 32

/* PAT9_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_OFFSET 16'h1634
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT9_EXE_CFG_INNER_WIDTH 32

/* PAT10_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_OFFSET 16'h1638
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT10_EXE_CFG_INNER_WIDTH 32

/* PAT11_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_OFFSET 16'h163c
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT11_EXE_CFG_INNER_WIDTH 32

/* PAT12_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_OFFSET 16'h1640
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT12_EXE_CFG_INNER_WIDTH 32

/* PAT13_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_OFFSET 16'h1644
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT13_EXE_CFG_INNER_WIDTH 32

/* PAT14_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_OFFSET 16'h1648
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT14_EXE_CFG_INNER_WIDTH 32

/* PAT15_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_OFFSET 16'h164c
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT15_EXE_CFG_INNER_WIDTH 32

/* PAT16_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_OFFSET 16'h1650
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT16_EXE_CFG_INNER_WIDTH 32

/* PAT17_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_OFFSET 16'h1654
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT17_EXE_CFG_INNER_WIDTH 32

/* PAT18_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_OFFSET 16'h1658
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT18_EXE_CFG_INNER_WIDTH 32

/* PAT19_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_OFFSET 16'h165c
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT19_EXE_CFG_INNER_WIDTH 32

/* PAT20_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_OFFSET 16'h1660
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT20_EXE_CFG_INNER_WIDTH 32

/* PAT21_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_OFFSET 16'h1664
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT21_EXE_CFG_INNER_WIDTH 32

/* PAT22_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_OFFSET 16'h1668
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT22_EXE_CFG_INNER_WIDTH 32

/* PAT23_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_OFFSET 16'h166c
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT23_EXE_CFG_INNER_WIDTH 32

/* PAT24_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_OFFSET 16'h1670
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT24_EXE_CFG_INNER_WIDTH 32

/* PAT25_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_OFFSET 16'h1674
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT25_EXE_CFG_INNER_WIDTH 32

/* PAT26_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_OFFSET 16'h1678
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT26_EXE_CFG_INNER_WIDTH 32

/* PAT27_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_OFFSET 16'h167c
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT27_EXE_CFG_INNER_WIDTH 32

/* PAT28_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_OFFSET 16'h1680
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT28_EXE_CFG_INNER_WIDTH 32

/* PAT29_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_OFFSET 16'h1684
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT29_EXE_CFG_INNER_WIDTH 32

/* PAT30_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_OFFSET 16'h1688
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT30_EXE_CFG_INNER_WIDTH 32

/* PAT31_EXE_CFG_INNER */
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_OFFSET 16'h168c
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_LOOP_DLY 8:0
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_LOOP_DLY_WIDTH 9
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_LOOP_CNT 14:9
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_LOOP_CNT_WIDTH 6
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_KEEP_PAT 15
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_KEEP_CAS 16
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_NXT_PAT_DLY 26:17
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_NXT_PAT_DLY_WIDTH 10
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT31_EXE_CFG_INNER_WIDTH 32

/* DEFAULT_PAT_EXE_CFG_OUTER */
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_OFFSET 16'h1690
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_DEFAULT_PAT_EXE_CFG_OUTER_WIDTH 32

/* PAT0_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_OFFSET 16'h1694
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT0_EXE_CFG_OUTER_WIDTH 32

/* PAT1_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_OFFSET 16'h1698
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT1_EXE_CFG_OUTER_WIDTH 32

/* PAT2_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_OFFSET 16'h169c
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT2_EXE_CFG_OUTER_WIDTH 32

/* PAT3_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_OFFSET 16'h16a0
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT3_EXE_CFG_OUTER_WIDTH 32

/* PAT4_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_OFFSET 16'h16a4
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT4_EXE_CFG_OUTER_WIDTH 32

/* PAT5_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_OFFSET 16'h16a8
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT5_EXE_CFG_OUTER_WIDTH 32

/* PAT6_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_OFFSET 16'h16ac
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT6_EXE_CFG_OUTER_WIDTH 32

/* PAT7_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_OFFSET 16'h16b0
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT7_EXE_CFG_OUTER_WIDTH 32

/* PAT8_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_OFFSET 16'h16b4
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT8_EXE_CFG_OUTER_WIDTH 32

/* PAT9_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_OFFSET 16'h16b8
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT9_EXE_CFG_OUTER_WIDTH 32

/* PAT10_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_OFFSET 16'h16bc
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT10_EXE_CFG_OUTER_WIDTH 32

/* PAT11_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_OFFSET 16'h16c0
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT11_EXE_CFG_OUTER_WIDTH 32

/* PAT12_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_OFFSET 16'h16c4
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT12_EXE_CFG_OUTER_WIDTH 32

/* PAT13_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_OFFSET 16'h16c8
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT13_EXE_CFG_OUTER_WIDTH 32

/* PAT14_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_OFFSET 16'h16cc
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT14_EXE_CFG_OUTER_WIDTH 32

/* PAT15_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_OFFSET 16'h16d0
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT15_EXE_CFG_OUTER_WIDTH 32

/* PAT16_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_OFFSET 16'h16d4
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT16_EXE_CFG_OUTER_WIDTH 32

/* PAT17_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_OFFSET 16'h16d8
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT17_EXE_CFG_OUTER_WIDTH 32

/* PAT18_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_OFFSET 16'h16dc
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT18_EXE_CFG_OUTER_WIDTH 32

/* PAT19_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_OFFSET 16'h16e0
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT19_EXE_CFG_OUTER_WIDTH 32

/* PAT20_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_OFFSET 16'h16e4
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT20_EXE_CFG_OUTER_WIDTH 32

/* PAT21_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_OFFSET 16'h16e8
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT21_EXE_CFG_OUTER_WIDTH 32

/* PAT22_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_OFFSET 16'h16ec
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT22_EXE_CFG_OUTER_WIDTH 32

/* PAT23_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_OFFSET 16'h16f0
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT23_EXE_CFG_OUTER_WIDTH 32

/* PAT24_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_OFFSET 16'h16f4
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT24_EXE_CFG_OUTER_WIDTH 32

/* PAT25_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_OFFSET 16'h16f8
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT25_EXE_CFG_OUTER_WIDTH 32

/* PAT26_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_OFFSET 16'h16fc
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT26_EXE_CFG_OUTER_WIDTH 32

/* PAT27_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_OFFSET 16'h1700
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT27_EXE_CFG_OUTER_WIDTH 32

/* PAT28_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_OFFSET 16'h1704
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT28_EXE_CFG_OUTER_WIDTH 32

/* PAT29_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_OFFSET 16'h1708
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT29_EXE_CFG_OUTER_WIDTH 32

/* PAT30_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_OFFSET 16'h170c
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT30_EXE_CFG_OUTER_WIDTH 32

/* PAT31_EXE_CFG_OUTER */
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_OFFSET 16'h1710
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_LOOP_CNT 9:0
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_LOOP_CNT_WIDTH 10
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_KEEP_PAT 10
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_KEEP_PAT_WIDTH 1
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_KEEP_CAS 11
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_KEEP_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_NXT_PAT_DLY 26:12
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_NXT_PAT_DLY_WIDTH 15
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_NXT_PAT_IDX 31:27
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_FLD_NXT_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT31_EXE_CFG_OUTER_WIDTH 32

/* PAT_EXE_CTRL */
`define DDRMC5_MAIN_PAT_EXE_CTRL_OFFSET 16'h1714
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_START 0
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_START_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_RST 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_RST_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_START_PAT_IDX 6:2
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_START_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_STOP_PAT_IDX 11:7
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_STOP_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK0 12
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK0_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK1 13
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK1_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK2 14
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK2_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK3 15
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CMD_ADDR_TCK3_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_DQ 16
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_DQ_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_DMDBI_DQS 17
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_DMDBI_DQS_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CAS 18
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_CAS_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LATCH_DEFAULT_PATTERN_EN 19
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LATCH_DEFAULT_PATTERN_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_INNER_CONFIG 20
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_INNER_CONFIG_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_OUTER_CONFIG 21
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_OUTER_CONFIG_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_PDA_DQ_MODE_EN 22
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_PDA_DQ_MODE_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_NIBBLE_WISE_DQ_EN 23
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_NIBBLE_WISE_DQ_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_STEPSIZE 24
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_LOAD_DEFAULT_STEPSIZE_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_RESERVED 31:25
`define DDRMC5_MAIN_PAT_EXE_CTRL_FLD_RESERVED_WIDTH 7
`define DDRMC5_MAIN_PAT_EXE_CTRL_WIDTH 25

/* PAT_DEFAULT_LOAD_ENABLE */
`define DDRMC5_MAIN_PAT_DEFAULT_LOAD_ENABLE_OFFSET 16'h1718
`define DDRMC5_MAIN_PAT_DEFAULT_LOAD_ENABLE_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT_DEFAULT_LOAD_ENABLE_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT_DEFAULT_LOAD_ENABLE_WIDTH 32

/* PAT_EXE_STATUS */
`define DDRMC5_MAIN_PAT_EXE_STATUS_OFFSET 16'h171c
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_DONE 0
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_DONE_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_BUSY 1
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_PAT_IDX 6:2
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_PAT_IDX_WIDTH 5
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_RESERVED 31:7
`define DDRMC5_MAIN_PAT_EXE_STATUS_FLD_RESERVED_WIDTH 25
`define DDRMC5_MAIN_PAT_EXE_STATUS_WIDTH 7

/* PAT_EXE2DATA_VLD_LATENCY */
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_OFFSET 16'h1720
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_LATENCY 7:0
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_LATENCY_WIDTH 8
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_EN 8
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_RESERVED 31:9
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_FLD_RESERVED_WIDTH 23
`define DDRMC5_MAIN_PAT_EXE2DATA_VLD_LATENCY_WIDTH 9

/* ED_DONE_STATUS_31_0 */
`define DDRMC5_MAIN_ED_DONE_STATUS_31_0_OFFSET 16'h1724
`define DDRMC5_MAIN_ED_DONE_STATUS_31_0_FLD_VAL 31:0
`define DDRMC5_MAIN_ED_DONE_STATUS_31_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ED_DONE_STATUS_31_0_WIDTH 32

/* ED_DONE_STATUS_63_32 */
`define DDRMC5_MAIN_ED_DONE_STATUS_63_32_OFFSET 16'h1728
`define DDRMC5_MAIN_ED_DONE_STATUS_63_32_FLD_VAL 31:0
`define DDRMC5_MAIN_ED_DONE_STATUS_63_32_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ED_DONE_STATUS_63_32_WIDTH 32

/* ED_DONE_STATUS_79_64 */
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_OFFSET 16'h172c
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_FLD_VAL 15:0
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ED_DONE_STATUS_79_64_WIDTH 16

/* ED_0_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_OFFSET 16'h1730
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_0_ITERATION_STATUS_WIDTH 18

/* ED_1_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_OFFSET 16'h1734
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_1_ITERATION_STATUS_WIDTH 18

/* ED_2_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_OFFSET 16'h1738
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_2_ITERATION_STATUS_WIDTH 18

/* ED_3_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_OFFSET 16'h173c
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_3_ITERATION_STATUS_WIDTH 18

/* ED_4_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_OFFSET 16'h1740
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_4_ITERATION_STATUS_WIDTH 18

/* ED_5_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_OFFSET 16'h1744
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_5_ITERATION_STATUS_WIDTH 18

/* ED_6_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_OFFSET 16'h1748
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_6_ITERATION_STATUS_WIDTH 18

/* ED_7_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_OFFSET 16'h174c
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_7_ITERATION_STATUS_WIDTH 18

/* ED_8_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_OFFSET 16'h1750
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_8_ITERATION_STATUS_WIDTH 18

/* ED_9_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_OFFSET 16'h1754
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_9_ITERATION_STATUS_WIDTH 18

/* ED_10_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_OFFSET 16'h1758
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_10_ITERATION_STATUS_WIDTH 18

/* ED_11_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_OFFSET 16'h175c
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_11_ITERATION_STATUS_WIDTH 18

/* ED_12_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_OFFSET 16'h1760
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_12_ITERATION_STATUS_WIDTH 18

/* ED_13_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_OFFSET 16'h1764
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_13_ITERATION_STATUS_WIDTH 18

/* ED_14_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_OFFSET 16'h1768
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_14_ITERATION_STATUS_WIDTH 18

/* ED_15_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_OFFSET 16'h176c
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_15_ITERATION_STATUS_WIDTH 18

/* ED_16_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_OFFSET 16'h1770
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_16_ITERATION_STATUS_WIDTH 18

/* ED_17_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_OFFSET 16'h1774
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_17_ITERATION_STATUS_WIDTH 18

/* ED_18_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_OFFSET 16'h1778
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_18_ITERATION_STATUS_WIDTH 18

/* ED_19_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_OFFSET 16'h177c
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_19_ITERATION_STATUS_WIDTH 18

/* ED_20_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_OFFSET 16'h1780
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_20_ITERATION_STATUS_WIDTH 18

/* ED_21_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_OFFSET 16'h1784
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_21_ITERATION_STATUS_WIDTH 18

/* ED_22_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_OFFSET 16'h1788
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_22_ITERATION_STATUS_WIDTH 18

/* ED_23_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_OFFSET 16'h178c
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_23_ITERATION_STATUS_WIDTH 18

/* ED_24_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_OFFSET 16'h1790
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_24_ITERATION_STATUS_WIDTH 18

/* ED_25_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_OFFSET 16'h1794
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_25_ITERATION_STATUS_WIDTH 18

/* ED_26_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_OFFSET 16'h1798
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_26_ITERATION_STATUS_WIDTH 18

/* ED_27_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_OFFSET 16'h179c
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_27_ITERATION_STATUS_WIDTH 18

/* ED_28_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_OFFSET 16'h17a0
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_28_ITERATION_STATUS_WIDTH 18

/* ED_29_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_OFFSET 16'h17a4
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_29_ITERATION_STATUS_WIDTH 18

/* ED_30_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_OFFSET 16'h17a8
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_30_ITERATION_STATUS_WIDTH 18

/* ED_31_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_OFFSET 16'h17ac
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_31_ITERATION_STATUS_WIDTH 18

/* ED_32_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_OFFSET 16'h17b0
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_32_ITERATION_STATUS_WIDTH 18

/* ED_33_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_OFFSET 16'h17b4
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_33_ITERATION_STATUS_WIDTH 18

/* ED_34_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_OFFSET 16'h17b8
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_34_ITERATION_STATUS_WIDTH 18

/* ED_35_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_OFFSET 16'h17bc
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_35_ITERATION_STATUS_WIDTH 18

/* ED_36_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_OFFSET 16'h17c0
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_36_ITERATION_STATUS_WIDTH 18

/* ED_37_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_OFFSET 16'h17c4
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_37_ITERATION_STATUS_WIDTH 18

/* ED_38_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_OFFSET 16'h17c8
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_38_ITERATION_STATUS_WIDTH 18

/* ED_39_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_OFFSET 16'h17cc
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_39_ITERATION_STATUS_WIDTH 18

/* ED_40_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_OFFSET 16'h17d0
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_40_ITERATION_STATUS_WIDTH 18

/* ED_41_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_OFFSET 16'h17d4
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_41_ITERATION_STATUS_WIDTH 18

/* ED_42_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_OFFSET 16'h17d8
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_42_ITERATION_STATUS_WIDTH 18

/* ED_43_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_OFFSET 16'h17dc
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_43_ITERATION_STATUS_WIDTH 18

/* ED_44_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_OFFSET 16'h17e0
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_44_ITERATION_STATUS_WIDTH 18

/* ED_45_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_OFFSET 16'h17e4
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_45_ITERATION_STATUS_WIDTH 18

/* ED_46_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_OFFSET 16'h17e8
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_46_ITERATION_STATUS_WIDTH 18

/* ED_47_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_OFFSET 16'h17ec
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_47_ITERATION_STATUS_WIDTH 18

/* ED_48_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_OFFSET 16'h17f0
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_48_ITERATION_STATUS_WIDTH 18

/* ED_49_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_OFFSET 16'h17f4
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_49_ITERATION_STATUS_WIDTH 18

/* ED_50_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_OFFSET 16'h17f8
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_50_ITERATION_STATUS_WIDTH 18

/* ED_51_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_OFFSET 16'h17fc
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_51_ITERATION_STATUS_WIDTH 18

/* ED_52_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_OFFSET 16'h1800
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_52_ITERATION_STATUS_WIDTH 18

/* ED_53_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_OFFSET 16'h1804
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_53_ITERATION_STATUS_WIDTH 18

/* ED_54_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_OFFSET 16'h1808
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_54_ITERATION_STATUS_WIDTH 18

/* ED_55_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_OFFSET 16'h180c
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_55_ITERATION_STATUS_WIDTH 18

/* ED_56_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_OFFSET 16'h1810
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_56_ITERATION_STATUS_WIDTH 18

/* ED_57_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_OFFSET 16'h1814
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_57_ITERATION_STATUS_WIDTH 18

/* ED_58_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_OFFSET 16'h1818
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_58_ITERATION_STATUS_WIDTH 18

/* ED_59_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_OFFSET 16'h181c
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_59_ITERATION_STATUS_WIDTH 18

/* ED_60_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_OFFSET 16'h1820
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_60_ITERATION_STATUS_WIDTH 18

/* ED_61_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_OFFSET 16'h1824
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_61_ITERATION_STATUS_WIDTH 18

/* ED_62_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_OFFSET 16'h1828
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_62_ITERATION_STATUS_WIDTH 18

/* ED_63_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_OFFSET 16'h182c
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_63_ITERATION_STATUS_WIDTH 18

/* ED_64_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_OFFSET 16'h1830
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_64_ITERATION_STATUS_WIDTH 18

/* ED_65_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_OFFSET 16'h1834
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_65_ITERATION_STATUS_WIDTH 18

/* ED_66_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_OFFSET 16'h1838
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_66_ITERATION_STATUS_WIDTH 18

/* ED_67_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_OFFSET 16'h183c
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_67_ITERATION_STATUS_WIDTH 18

/* ED_68_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_OFFSET 16'h1840
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_68_ITERATION_STATUS_WIDTH 18

/* ED_69_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_OFFSET 16'h1844
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_69_ITERATION_STATUS_WIDTH 18

/* ED_70_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_OFFSET 16'h1848
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_70_ITERATION_STATUS_WIDTH 18

/* ED_71_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_OFFSET 16'h184c
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_71_ITERATION_STATUS_WIDTH 18

/* ED_72_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_OFFSET 16'h1850
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_72_ITERATION_STATUS_WIDTH 18

/* ED_73_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_OFFSET 16'h1854
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_73_ITERATION_STATUS_WIDTH 18

/* ED_74_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_OFFSET 16'h1858
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_74_ITERATION_STATUS_WIDTH 18

/* ED_75_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_OFFSET 16'h185c
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_75_ITERATION_STATUS_WIDTH 18

/* ED_76_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_OFFSET 16'h1860
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_76_ITERATION_STATUS_WIDTH 18

/* ED_77_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_OFFSET 16'h1864
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_77_ITERATION_STATUS_WIDTH 18

/* ED_78_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_OFFSET 16'h1868
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_78_ITERATION_STATUS_WIDTH 18

/* ED_79_ITERATION_STATUS */
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_OFFSET 16'h186c
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_ITR_COUNTS 8:0
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_ITR_COUNTS_WIDTH 9
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_LAST_VALID_WIN 17:9
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_LAST_VALID_WIN_WIDTH 9
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_RESERVED 31:18
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_FLD_RESERVED_WIDTH 14
`define DDRMC5_MAIN_ED_79_ITERATION_STATUS_WIDTH 18

/* ED_CONFIG */
`define DDRMC5_MAIN_ED_CONFIG_OFFSET 16'h1870
`define DDRMC5_MAIN_ED_CONFIG_FLD_RST 0
`define DDRMC5_MAIN_ED_CONFIG_FLD_RST_WIDTH 1
`define DDRMC5_MAIN_ED_CONFIG_FLD_SET1 1
`define DDRMC5_MAIN_ED_CONFIG_FLD_SET1_WIDTH 1
`define DDRMC5_MAIN_ED_CONFIG_FLD_SET0 2
`define DDRMC5_MAIN_ED_CONFIG_FLD_SET0_WIDTH 1
`define DDRMC5_MAIN_ED_CONFIG_FLD_ANALYZE 3
`define DDRMC5_MAIN_ED_CONFIG_FLD_ANALYZE_WIDTH 1
`define DDRMC5_MAIN_ED_CONFIG_FLD_MODE 5:4
`define DDRMC5_MAIN_ED_CONFIG_FLD_MODE_WIDTH 2
`define DDRMC5_MAIN_ED_CONFIG_FLD_MIN_VALID_WIN 13:6
`define DDRMC5_MAIN_ED_CONFIG_FLD_MIN_VALID_WIN_WIDTH 8
`define DDRMC5_MAIN_ED_CONFIG_FLD_RESERVED 31:14
`define DDRMC5_MAIN_ED_CONFIG_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_ED_CONFIG_WIDTH 14

/* ED_31_0_MASK */
`define DDRMC5_MAIN_ED_31_0_MASK_OFFSET 16'h1874
`define DDRMC5_MAIN_ED_31_0_MASK_FLD_VAL 31:0
`define DDRMC5_MAIN_ED_31_0_MASK_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ED_31_0_MASK_WIDTH 32

/* ED_63_32_MASK */
`define DDRMC5_MAIN_ED_63_32_MASK_OFFSET 16'h1878
`define DDRMC5_MAIN_ED_63_32_MASK_FLD_VAL 31:0
`define DDRMC5_MAIN_ED_63_32_MASK_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ED_63_32_MASK_WIDTH 32

/* ED_79_64_MASK */
`define DDRMC5_MAIN_ED_79_64_MASK_OFFSET 16'h187c
`define DDRMC5_MAIN_ED_79_64_MASK_FLD_VAL 15:0
`define DDRMC5_MAIN_ED_79_64_MASK_FLD_VAL_WIDTH 16
`define DDRMC5_MAIN_ED_79_64_MASK_FLD_RESERVED 31:16
`define DDRMC5_MAIN_ED_79_64_MASK_FLD_RESERVED_WIDTH 16
`define DDRMC5_MAIN_ED_79_64_MASK_WIDTH 16

/* CMP2ED_STATUS_CONFIG */
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_OFFSET 16'h1880
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_CMP_TYPE 2:0
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_CMP_TYPE_WIDTH 3
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_CMP_EDGE 5:3
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_CMP_EDGE_WIDTH 3
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_RESERVED 31:6
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_FLD_RESERVED_WIDTH 26
`define DDRMC5_MAIN_CMP2ED_STATUS_CONFIG_WIDTH 6

/* ACC_CTRL */
`define DDRMC5_MAIN_ACC_CTRL_OFFSET 16'h1884
`define DDRMC5_MAIN_ACC_CTRL_FLD_START 0
`define DDRMC5_MAIN_ACC_CTRL_FLD_START_WIDTH 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_RST 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_RST_WIDTH 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_STOP 2
`define DDRMC5_MAIN_ACC_CTRL_FLD_STOP_WIDTH 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_TIMER_STOP 3
`define DDRMC5_MAIN_ACC_CTRL_FLD_TIMER_STOP_WIDTH 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_WCMPR_CLR 4
`define DDRMC5_MAIN_ACC_CTRL_FLD_WCMPR_CLR_WIDTH 1
`define DDRMC5_MAIN_ACC_CTRL_FLD_PATTERN_GEN_MODE 7:5
`define DDRMC5_MAIN_ACC_CTRL_FLD_PATTERN_GEN_MODE_WIDTH 3
`define DDRMC5_MAIN_ACC_CTRL_FLD_RESERVED 31:8
`define DDRMC5_MAIN_ACC_CTRL_FLD_RESERVED_WIDTH 24
`define DDRMC5_MAIN_ACC_CTRL_WIDTH 8

/* ACC_STATUS */
`define DDRMC5_MAIN_ACC_STATUS_OFFSET 16'h1888
`define DDRMC5_MAIN_ACC_STATUS_FLD_DONE 0
`define DDRMC5_MAIN_ACC_STATUS_FLD_DONE_WIDTH 1
`define DDRMC5_MAIN_ACC_STATUS_FLD_BUSY 1
`define DDRMC5_MAIN_ACC_STATUS_FLD_BUSY_WIDTH 1
`define DDRMC5_MAIN_ACC_STATUS_FLD_ERROR 2
`define DDRMC5_MAIN_ACC_STATUS_FLD_ERROR_WIDTH 1
`define DDRMC5_MAIN_ACC_STATUS_FLD_STAGE 6:3
`define DDRMC5_MAIN_ACC_STATUS_FLD_STAGE_WIDTH 4
`define DDRMC5_MAIN_ACC_STATUS_FLD_ITERATION 16:7
`define DDRMC5_MAIN_ACC_STATUS_FLD_ITERATION_WIDTH 10
`define DDRMC5_MAIN_ACC_STATUS_FLD_RESERVED 31:17
`define DDRMC5_MAIN_ACC_STATUS_FLD_RESERVED_WIDTH 15
`define DDRMC5_MAIN_ACC_STATUS_WIDTH 17

/* ACC_PAT_WAIT_LIMIT */
`define DDRMC5_MAIN_ACC_PAT_WAIT_LIMIT_OFFSET 16'h188c
`define DDRMC5_MAIN_ACC_PAT_WAIT_LIMIT_FLD_VAL 31:0
`define DDRMC5_MAIN_ACC_PAT_WAIT_LIMIT_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ACC_PAT_WAIT_LIMIT_WIDTH 32

/* ACC_RPI_WAIT_LIMIT */
`define DDRMC5_MAIN_ACC_RPI_WAIT_LIMIT_OFFSET 16'h1890
`define DDRMC5_MAIN_ACC_RPI_WAIT_LIMIT_FLD_VAL 31:0
`define DDRMC5_MAIN_ACC_RPI_WAIT_LIMIT_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ACC_RPI_WAIT_LIMIT_WIDTH 32

/* ACC_ITR_LIMIT */
`define DDRMC5_MAIN_ACC_ITR_LIMIT_OFFSET 16'h1894
`define DDRMC5_MAIN_ACC_ITR_LIMIT_FLD_VAL 31:0
`define DDRMC5_MAIN_ACC_ITR_LIMIT_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ACC_ITR_LIMIT_WIDTH 32

/* PAT_END2ED_EN_DELAY */
`define DDRMC5_MAIN_PAT_END2ED_EN_DELAY_OFFSET 16'h1898
`define DDRMC5_MAIN_PAT_END2ED_EN_DELAY_FLD_VAL 31:0
`define DDRMC5_MAIN_PAT_END2ED_EN_DELAY_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_PAT_END2ED_EN_DELAY_WIDTH 32

/* ACC_PAT_START_DELAY */
`define DDRMC5_MAIN_ACC_PAT_START_DELAY_OFFSET 16'h189c
`define DDRMC5_MAIN_ACC_PAT_START_DELAY_FLD_VAL 31:0
`define DDRMC5_MAIN_ACC_PAT_START_DELAY_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_ACC_PAT_START_DELAY_WIDTH 32

/* POST_DELAY_UPDATE_DELAY */
`define DDRMC5_MAIN_POST_DELAY_UPDATE_DELAY_OFFSET 16'h18a0
`define DDRMC5_MAIN_POST_DELAY_UPDATE_DELAY_FLD_VAL 31:0
`define DDRMC5_MAIN_POST_DELAY_UPDATE_DELAY_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_POST_DELAY_UPDATE_DELAY_WIDTH 32

/* PAT_LOW_FEQ_MODE */
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_OFFSET 16'h18a4
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_FLD_EN 0
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_FLD_RESERVED 31:1
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_PAT_LOW_FEQ_MODE_WIDTH 1

/* CAL_DEBUG_REG_0 */
`define DDRMC5_MAIN_CAL_DEBUG_REG_0_OFFSET 16'h18a8
`define DDRMC5_MAIN_CAL_DEBUG_REG_0_FLD_VAL 31:0
`define DDRMC5_MAIN_CAL_DEBUG_REG_0_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_CAL_DEBUG_REG_0_WIDTH 32

/* CAL_DEBUG_REG_1 */
`define DDRMC5_MAIN_CAL_DEBUG_REG_1_OFFSET 16'h18ac
`define DDRMC5_MAIN_CAL_DEBUG_REG_1_FLD_VAL 31:0
`define DDRMC5_MAIN_CAL_DEBUG_REG_1_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_CAL_DEBUG_REG_1_WIDTH 32

/* CAL_DEBUG_REG_2 */
`define DDRMC5_MAIN_CAL_DEBUG_REG_2_OFFSET 16'h18b0
`define DDRMC5_MAIN_CAL_DEBUG_REG_2_FLD_VAL 31:0
`define DDRMC5_MAIN_CAL_DEBUG_REG_2_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_CAL_DEBUG_REG_2_WIDTH 32

/* CAL_DEBUG_REG_3 */
`define DDRMC5_MAIN_CAL_DEBUG_REG_3_OFFSET 16'h18b4
`define DDRMC5_MAIN_CAL_DEBUG_REG_3_FLD_VAL 31:0
`define DDRMC5_MAIN_CAL_DEBUG_REG_3_FLD_VAL_WIDTH 32
`define DDRMC5_MAIN_CAL_DEBUG_REG_3_WIDTH 32

/* XPI_DQS_CNTRL */
`define DDRMC5_MAIN_XPI_DQS_CNTRL_OFFSET 16'h18b8
`define DDRMC5_MAIN_XPI_DQS_CNTRL_FLD_EN 0
`define DDRMC5_MAIN_XPI_DQS_CNTRL_FLD_EN_WIDTH 1
`define DDRMC5_MAIN_XPI_DQS_CNTRL_FLD_RESERVED 31:1
`define DDRMC5_MAIN_XPI_DQS_CNTRL_FLD_RESERVED_WIDTH 31
`define DDRMC5_MAIN_XPI_DQS_CNTRL_WIDTH 1

/* PAT0_STEPSIZE */
`define DDRMC5_MAIN_PAT0_STEPSIZE_OFFSET 16'h18bc
`define DDRMC5_MAIN_PAT0_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT0_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT0_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT0_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT0_STEPSIZE_WIDTH 14

/* PAT1_STEPSIZE */
`define DDRMC5_MAIN_PAT1_STEPSIZE_OFFSET 16'h18c0
`define DDRMC5_MAIN_PAT1_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT1_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT1_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT1_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT1_STEPSIZE_WIDTH 14

/* PAT2_STEPSIZE */
`define DDRMC5_MAIN_PAT2_STEPSIZE_OFFSET 16'h18c4
`define DDRMC5_MAIN_PAT2_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT2_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT2_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT2_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT2_STEPSIZE_WIDTH 14

/* PAT3_STEPSIZE */
`define DDRMC5_MAIN_PAT3_STEPSIZE_OFFSET 16'h18c8
`define DDRMC5_MAIN_PAT3_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT3_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT3_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT3_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT3_STEPSIZE_WIDTH 14

/* PAT4_STEPSIZE */
`define DDRMC5_MAIN_PAT4_STEPSIZE_OFFSET 16'h18cc
`define DDRMC5_MAIN_PAT4_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT4_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT4_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT4_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT4_STEPSIZE_WIDTH 14

/* PAT5_STEPSIZE */
`define DDRMC5_MAIN_PAT5_STEPSIZE_OFFSET 16'h18d0
`define DDRMC5_MAIN_PAT5_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT5_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT5_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT5_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT5_STEPSIZE_WIDTH 14

/* PAT6_STEPSIZE */
`define DDRMC5_MAIN_PAT6_STEPSIZE_OFFSET 16'h18d4
`define DDRMC5_MAIN_PAT6_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT6_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT6_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT6_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT6_STEPSIZE_WIDTH 14

/* PAT7_STEPSIZE */
`define DDRMC5_MAIN_PAT7_STEPSIZE_OFFSET 16'h18d8
`define DDRMC5_MAIN_PAT7_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT7_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT7_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT7_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT7_STEPSIZE_WIDTH 14

/* PAT8_STEPSIZE */
`define DDRMC5_MAIN_PAT8_STEPSIZE_OFFSET 16'h18dc
`define DDRMC5_MAIN_PAT8_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT8_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT8_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT8_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT8_STEPSIZE_WIDTH 14

/* PAT9_STEPSIZE */
`define DDRMC5_MAIN_PAT9_STEPSIZE_OFFSET 16'h18e0
`define DDRMC5_MAIN_PAT9_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT9_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT9_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT9_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT9_STEPSIZE_WIDTH 14

/* PAT10_STEPSIZE */
`define DDRMC5_MAIN_PAT10_STEPSIZE_OFFSET 16'h18e4
`define DDRMC5_MAIN_PAT10_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT10_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT10_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT10_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT10_STEPSIZE_WIDTH 14

/* PAT11_STEPSIZE */
`define DDRMC5_MAIN_PAT11_STEPSIZE_OFFSET 16'h18e8
`define DDRMC5_MAIN_PAT11_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT11_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT11_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT11_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT11_STEPSIZE_WIDTH 14

/* PAT12_STEPSIZE */
`define DDRMC5_MAIN_PAT12_STEPSIZE_OFFSET 16'h18ec
`define DDRMC5_MAIN_PAT12_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT12_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT12_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT12_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT12_STEPSIZE_WIDTH 14

/* PAT13_STEPSIZE */
`define DDRMC5_MAIN_PAT13_STEPSIZE_OFFSET 16'h18f0
`define DDRMC5_MAIN_PAT13_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT13_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT13_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT13_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT13_STEPSIZE_WIDTH 14

/* PAT14_STEPSIZE */
`define DDRMC5_MAIN_PAT14_STEPSIZE_OFFSET 16'h18f4
`define DDRMC5_MAIN_PAT14_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT14_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT14_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT14_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT14_STEPSIZE_WIDTH 14

/* PAT15_STEPSIZE */
`define DDRMC5_MAIN_PAT15_STEPSIZE_OFFSET 16'h18f8
`define DDRMC5_MAIN_PAT15_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT15_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT15_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT15_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT15_STEPSIZE_WIDTH 14

/* PAT16_STEPSIZE */
`define DDRMC5_MAIN_PAT16_STEPSIZE_OFFSET 16'h18fc
`define DDRMC5_MAIN_PAT16_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT16_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT16_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT16_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT16_STEPSIZE_WIDTH 14

/* PAT17_STEPSIZE */
`define DDRMC5_MAIN_PAT17_STEPSIZE_OFFSET 16'h1900
`define DDRMC5_MAIN_PAT17_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT17_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT17_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT17_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT17_STEPSIZE_WIDTH 14

/* PAT18_STEPSIZE */
`define DDRMC5_MAIN_PAT18_STEPSIZE_OFFSET 16'h1904
`define DDRMC5_MAIN_PAT18_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT18_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT18_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT18_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT18_STEPSIZE_WIDTH 14

/* PAT19_STEPSIZE */
`define DDRMC5_MAIN_PAT19_STEPSIZE_OFFSET 16'h1908
`define DDRMC5_MAIN_PAT19_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT19_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT19_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT19_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT19_STEPSIZE_WIDTH 14

/* PAT20_STEPSIZE */
`define DDRMC5_MAIN_PAT20_STEPSIZE_OFFSET 16'h190c
`define DDRMC5_MAIN_PAT20_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT20_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT20_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT20_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT20_STEPSIZE_WIDTH 14

/* PAT21_STEPSIZE */
`define DDRMC5_MAIN_PAT21_STEPSIZE_OFFSET 16'h1910
`define DDRMC5_MAIN_PAT21_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT21_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT21_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT21_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT21_STEPSIZE_WIDTH 14

/* PAT22_STEPSIZE */
`define DDRMC5_MAIN_PAT22_STEPSIZE_OFFSET 16'h1914
`define DDRMC5_MAIN_PAT22_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT22_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT22_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT22_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT22_STEPSIZE_WIDTH 14

/* PAT23_STEPSIZE */
`define DDRMC5_MAIN_PAT23_STEPSIZE_OFFSET 16'h1918
`define DDRMC5_MAIN_PAT23_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT23_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT23_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT23_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT23_STEPSIZE_WIDTH 14

/* PAT24_STEPSIZE */
`define DDRMC5_MAIN_PAT24_STEPSIZE_OFFSET 16'h191c
`define DDRMC5_MAIN_PAT24_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT24_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT24_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT24_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT24_STEPSIZE_WIDTH 14

/* PAT25_STEPSIZE */
`define DDRMC5_MAIN_PAT25_STEPSIZE_OFFSET 16'h1920
`define DDRMC5_MAIN_PAT25_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT25_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT25_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT25_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT25_STEPSIZE_WIDTH 14

/* PAT26_STEPSIZE */
`define DDRMC5_MAIN_PAT26_STEPSIZE_OFFSET 16'h1924
`define DDRMC5_MAIN_PAT26_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT26_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT26_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT26_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT26_STEPSIZE_WIDTH 14

/* PAT27_STEPSIZE */
`define DDRMC5_MAIN_PAT27_STEPSIZE_OFFSET 16'h1928
`define DDRMC5_MAIN_PAT27_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT27_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT27_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT27_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT27_STEPSIZE_WIDTH 14

/* PAT28_STEPSIZE */
`define DDRMC5_MAIN_PAT28_STEPSIZE_OFFSET 16'h192c
`define DDRMC5_MAIN_PAT28_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT28_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT28_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT28_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT28_STEPSIZE_WIDTH 14

/* PAT29_STEPSIZE */
`define DDRMC5_MAIN_PAT29_STEPSIZE_OFFSET 16'h1930
`define DDRMC5_MAIN_PAT29_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT29_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT29_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT29_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT29_STEPSIZE_WIDTH 14

/* PAT30_STEPSIZE */
`define DDRMC5_MAIN_PAT30_STEPSIZE_OFFSET 16'h1934
`define DDRMC5_MAIN_PAT30_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT30_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT30_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT30_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT30_STEPSIZE_WIDTH 14

/* PAT31_STEPSIZE */
`define DDRMC5_MAIN_PAT31_STEPSIZE_OFFSET 16'h1938
`define DDRMC5_MAIN_PAT31_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT31_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT31_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT31_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT31_STEPSIZE_WIDTH 14

/* PAT_DEFAULT_STEPSIZE */
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_OFFSET 16'h193c
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_FLD_VAL 13:0
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_FLD_VAL_WIDTH 14
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_FLD_RESERVED 31:14
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_FLD_RESERVED_WIDTH 18
`define DDRMC5_MAIN_PAT_DEFAULT_STEPSIZE_WIDTH 14

/* DDR5_SPARE_STAT_CFG0 */
`define DDRMC5_MAIN_DDR5_SPARE_STAT_CFG0_OFFSET 16'h1940
`define DDRMC5_MAIN_DDR5_SPARE_STAT_CFG0_FLD_SPARE 31:0
`define DDRMC5_MAIN_DDR5_SPARE_STAT_CFG0_FLD_SPARE_WIDTH 32
`define DDRMC5_MAIN_DDR5_SPARE_STAT_CFG0_WIDTH 32

// spyglass enable_block ConstName
`endif
