module matvec (
		input  wire        clock,  //  clock.clk
		input  wire        resetn, //  reset.reset_n
		input  wire        start,  //   call.valid
		output wire        busy,   //       .stall
		output wire        done,   // return.valid
		input  wire        stall,  //       .stall
		input  wire [63:0] M,      //      M.data
		input  wire [63:0] V,      //      V.data
		input  wire [63:0] Out0    //   Out0.data
	);
endmodule

