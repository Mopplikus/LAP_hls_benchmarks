// jacobi_1d.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module jacobi_1d (
		input  wire        clock,  //  clock.clk
		input  wire        resetn, //  reset.reset_n
		input  wire        start,  //   call.valid
		output wire        busy,   //       .stall
		output wire        done,   // return.valid
		input  wire        stall,  //       .stall
		input  wire [63:0] A_1,    //    A_1.data
		input  wire [63:0] A_2,    //    A_2.data
		input  wire [63:0] B       //      B.data
	);

	jacobi_1d_internal jacobi_1d_internal_inst (
		.clock  (clock),  //   input,   width = 1,  clock.clk
		.resetn (resetn), //   input,   width = 1,  reset.reset_n
		.start  (start),  //   input,   width = 1,   call.valid
		.busy   (busy),   //  output,   width = 1,       .stall
		.done   (done),   //  output,   width = 1, return.valid
		.stall  (stall),  //   input,   width = 1,       .stall
		.A_1    (A_1),    //   input,  width = 64,    A_1.data
		.A_2    (A_2),    //   input,  width = 64,    A_2.data
		.B      (B)       //   input,  width = 64,      B.data
	);

endmodule
