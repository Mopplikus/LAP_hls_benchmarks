`ifndef BFM_SIMULATION
`define EN_XPI_IF
`endif
`include "noc_define.vh"
`include "noc2_npp_ddrmc5_define.vh"
`include "noc_ddrmc5_define.vh"
`include "noc_npp_common_define.vh"
`include "ddr5mc_na_common_define.vh"
`include "ddr5mc_dc_common_define.vh"
`include "ddr5mc_bfm_na_noc_regs_defines.vh"
`include "ddr5mc_bfm_main_regs_defines.vh"
`include "ddr5mc_bfm_macros.svh"
`include "ddr5mc_bfm_top_io_define.vh"
`include "ddr5mc_bfm_cal_common_define.vh"
