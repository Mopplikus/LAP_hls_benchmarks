	component if_loop_3 is
		port (
			clock      : in  std_logic                     := 'X';             -- clk
			resetn     : in  std_logic                     := 'X';             -- reset_n
			start      : in  std_logic                     := 'X';             -- valid
			busy       : out std_logic;                                        -- stall
			done       : out std_logic;                                        -- valid
			stall      : in  std_logic                     := 'X';             -- stall
			returndata : out std_logic_vector(31 downto 0);                    -- data
			a          : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			b          : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			n          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- data
		);
	end component if_loop_3;

	u0 : component if_loop_3
		port map (
			clock      => CONNECTED_TO_clock,      --      clock.clk
			resetn     => CONNECTED_TO_resetn,     --      reset.reset_n
			start      => CONNECTED_TO_start,      --       call.valid
			busy       => CONNECTED_TO_busy,       --           .stall
			done       => CONNECTED_TO_done,       --     return.valid
			stall      => CONNECTED_TO_stall,      --           .stall
			returndata => CONNECTED_TO_returndata, -- returndata.data
			a          => CONNECTED_TO_a,          --          a.data
			b          => CONNECTED_TO_b,          --          b.data
			n          => CONNECTED_TO_n           --          n.data
		);

