module STORE_QUEUE_LSQ_E( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_8, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_9, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_10, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_11, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_12, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_13, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_14, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_15, // @[:@6.4]
  input         io_bbStorePorts_0, // @[:@6.4]
  input         io_bbNumStores, // @[:@6.4]
  output [3:0]  io_storeTail, // @[:@6.4]
  output [3:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [3:0]  io_loadTail, // @[:@6.4]
  input  [3:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadAddressDone_8, // @[:@6.4]
  input         io_loadAddressDone_9, // @[:@6.4]
  input         io_loadAddressDone_10, // @[:@6.4]
  input         io_loadAddressDone_11, // @[:@6.4]
  input         io_loadAddressDone_12, // @[:@6.4]
  input         io_loadAddressDone_13, // @[:@6.4]
  input         io_loadAddressDone_14, // @[:@6.4]
  input         io_loadAddressDone_15, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input         io_loadDataDone_8, // @[:@6.4]
  input         io_loadDataDone_9, // @[:@6.4]
  input         io_loadDataDone_10, // @[:@6.4]
  input         io_loadDataDone_11, // @[:@6.4]
  input         io_loadDataDone_12, // @[:@6.4]
  input         io_loadDataDone_13, // @[:@6.4]
  input         io_loadDataDone_14, // @[:@6.4]
  input         io_loadDataDone_15, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_7, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_8, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_9, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_10, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_11, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_12, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_13, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_14, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_15, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeAddrDone_8, // @[:@6.4]
  output        io_storeAddrDone_9, // @[:@6.4]
  output        io_storeAddrDone_10, // @[:@6.4]
  output        io_storeAddrDone_11, // @[:@6.4]
  output        io_storeAddrDone_12, // @[:@6.4]
  output        io_storeAddrDone_13, // @[:@6.4]
  output        io_storeAddrDone_14, // @[:@6.4]
  output        io_storeAddrDone_15, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output        io_storeDataDone_8, // @[:@6.4]
  output        io_storeDataDone_9, // @[:@6.4]
  output        io_storeDataDone_10, // @[:@6.4]
  output        io_storeDataDone_11, // @[:@6.4]
  output        io_storeDataDone_12, // @[:@6.4]
  output        io_storeDataDone_13, // @[:@6.4]
  output        io_storeDataDone_14, // @[:@6.4]
  output        io_storeDataDone_15, // @[:@6.4]
  output [31:0] io_storeAddrQueue_0, // @[:@6.4]
  output [31:0] io_storeAddrQueue_1, // @[:@6.4]
  output [31:0] io_storeAddrQueue_2, // @[:@6.4]
  output [31:0] io_storeAddrQueue_3, // @[:@6.4]
  output [31:0] io_storeAddrQueue_4, // @[:@6.4]
  output [31:0] io_storeAddrQueue_5, // @[:@6.4]
  output [31:0] io_storeAddrQueue_6, // @[:@6.4]
  output [31:0] io_storeAddrQueue_7, // @[:@6.4]
  output [31:0] io_storeAddrQueue_8, // @[:@6.4]
  output [31:0] io_storeAddrQueue_9, // @[:@6.4]
  output [31:0] io_storeAddrQueue_10, // @[:@6.4]
  output [31:0] io_storeAddrQueue_11, // @[:@6.4]
  output [31:0] io_storeAddrQueue_12, // @[:@6.4]
  output [31:0] io_storeAddrQueue_13, // @[:@6.4]
  output [31:0] io_storeAddrQueue_14, // @[:@6.4]
  output [31:0] io_storeAddrQueue_15, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_8, // @[:@6.4]
  output [31:0] io_storeDataQueue_9, // @[:@6.4]
  output [31:0] io_storeDataQueue_10, // @[:@6.4]
  output [31:0] io_storeDataQueue_11, // @[:@6.4]
  output [31:0] io_storeDataQueue_12, // @[:@6.4]
  output [31:0] io_storeDataQueue_13, // @[:@6.4]
  output [31:0] io_storeDataQueue_14, // @[:@6.4]
  output [31:0] io_storeDataQueue_15, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input         io_storeDataEnable_1, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_1, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input         io_storeAddrEnable_1, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_0, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_1, // @[:@6.4]
  output [31:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  output        io_storeEnableToMem, // @[:@6.4]
  input         io_memIsReadyForStores // @[:@6.4]
);
  reg [3:0] head; // @[StoreQueue.scala 50:21:@8.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[StoreQueue.scala 51:21:@9.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_97;
  reg  allocatedEntries_0; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_98;
  reg  allocatedEntries_1; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_99;
  reg  allocatedEntries_2; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_100;
  reg  allocatedEntries_3; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_101;
  reg  allocatedEntries_4; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_102;
  reg  allocatedEntries_5; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_103;
  reg  allocatedEntries_6; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_104;
  reg  allocatedEntries_7; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_105;
  reg  allocatedEntries_8; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_106;
  reg  allocatedEntries_9; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_107;
  reg  allocatedEntries_10; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_108;
  reg  allocatedEntries_11; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_109;
  reg  allocatedEntries_12; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_110;
  reg  allocatedEntries_13; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_111;
  reg  allocatedEntries_14; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_112;
  reg  allocatedEntries_15; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_113;
  reg  storeCompleted_0; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_114;
  reg  storeCompleted_1; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_115;
  reg  storeCompleted_2; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_116;
  reg  storeCompleted_3; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_117;
  reg  storeCompleted_4; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_118;
  reg  storeCompleted_5; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_119;
  reg  storeCompleted_6; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_120;
  reg  storeCompleted_7; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_121;
  reg  storeCompleted_8; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_122;
  reg  storeCompleted_9; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_123;
  reg  storeCompleted_10; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_124;
  reg  storeCompleted_11; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_125;
  reg  storeCompleted_12; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_126;
  reg  storeCompleted_13; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_127;
  reg  storeCompleted_14; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_128;
  reg  storeCompleted_15; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_129;
  reg  checkBits_0; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_130;
  reg  checkBits_1; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_131;
  reg  checkBits_2; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_132;
  reg  checkBits_3; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_133;
  reg  checkBits_4; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_134;
  reg  checkBits_5; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_135;
  reg  checkBits_6; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_136;
  reg  checkBits_7; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_137;
  reg  checkBits_8; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_138;
  reg  checkBits_9; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_139;
  reg  checkBits_10; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_140;
  reg  checkBits_11; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_141;
  reg  checkBits_12; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_142;
  reg  checkBits_13; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_143;
  reg  checkBits_14; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_144;
  reg  checkBits_15; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_145;
  wire [5:0] _GEN_1202; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1604; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1605; // @[util.scala 14:20:@174.4]
  wire [5:0] _T_1606; // @[util.scala 14:20:@175.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@176.4]
  wire [4:0] _T_1607; // @[util.scala 14:25:@176.4]
  wire [4:0] _GEN_1203; // @[StoreQueue.scala 70:46:@177.4]
  wire  _T_1608; // @[StoreQueue.scala 70:46:@177.4]
  wire  initBits_0; // @[StoreQueue.scala 70:64:@178.4]
  wire [6:0] _T_1613; // @[util.scala 14:20:@180.4]
  wire [6:0] _T_1614; // @[util.scala 14:20:@181.4]
  wire [5:0] _T_1615; // @[util.scala 14:20:@182.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@183.4]
  wire [4:0] _T_1616; // @[util.scala 14:25:@183.4]
  wire  _T_1617; // @[StoreQueue.scala 70:46:@184.4]
  wire  initBits_1; // @[StoreQueue.scala 70:64:@185.4]
  wire [6:0] _T_1622; // @[util.scala 14:20:@187.4]
  wire [6:0] _T_1623; // @[util.scala 14:20:@188.4]
  wire [5:0] _T_1624; // @[util.scala 14:20:@189.4]
  wire [5:0] _GEN_34; // @[util.scala 14:25:@190.4]
  wire [4:0] _T_1625; // @[util.scala 14:25:@190.4]
  wire  _T_1626; // @[StoreQueue.scala 70:46:@191.4]
  wire  initBits_2; // @[StoreQueue.scala 70:64:@192.4]
  wire [6:0] _T_1631; // @[util.scala 14:20:@194.4]
  wire [6:0] _T_1632; // @[util.scala 14:20:@195.4]
  wire [5:0] _T_1633; // @[util.scala 14:20:@196.4]
  wire [5:0] _GEN_50; // @[util.scala 14:25:@197.4]
  wire [4:0] _T_1634; // @[util.scala 14:25:@197.4]
  wire  _T_1635; // @[StoreQueue.scala 70:46:@198.4]
  wire  initBits_3; // @[StoreQueue.scala 70:64:@199.4]
  wire [6:0] _T_1640; // @[util.scala 14:20:@201.4]
  wire [6:0] _T_1641; // @[util.scala 14:20:@202.4]
  wire [5:0] _T_1642; // @[util.scala 14:20:@203.4]
  wire [5:0] _GEN_68; // @[util.scala 14:25:@204.4]
  wire [4:0] _T_1643; // @[util.scala 14:25:@204.4]
  wire  _T_1644; // @[StoreQueue.scala 70:46:@205.4]
  wire  initBits_4; // @[StoreQueue.scala 70:64:@206.4]
  wire [6:0] _T_1649; // @[util.scala 14:20:@208.4]
  wire [6:0] _T_1650; // @[util.scala 14:20:@209.4]
  wire [5:0] _T_1651; // @[util.scala 14:20:@210.4]
  wire [5:0] _GEN_84; // @[util.scala 14:25:@211.4]
  wire [4:0] _T_1652; // @[util.scala 14:25:@211.4]
  wire  _T_1653; // @[StoreQueue.scala 70:46:@212.4]
  wire  initBits_5; // @[StoreQueue.scala 70:64:@213.4]
  wire [6:0] _T_1658; // @[util.scala 14:20:@215.4]
  wire [6:0] _T_1659; // @[util.scala 14:20:@216.4]
  wire [5:0] _T_1660; // @[util.scala 14:20:@217.4]
  wire [5:0] _GEN_102; // @[util.scala 14:25:@218.4]
  wire [4:0] _T_1661; // @[util.scala 14:25:@218.4]
  wire  _T_1662; // @[StoreQueue.scala 70:46:@219.4]
  wire  initBits_6; // @[StoreQueue.scala 70:64:@220.4]
  wire [6:0] _T_1667; // @[util.scala 14:20:@222.4]
  wire [6:0] _T_1668; // @[util.scala 14:20:@223.4]
  wire [5:0] _T_1669; // @[util.scala 14:20:@224.4]
  wire [5:0] _GEN_118; // @[util.scala 14:25:@225.4]
  wire [4:0] _T_1670; // @[util.scala 14:25:@225.4]
  wire  _T_1671; // @[StoreQueue.scala 70:46:@226.4]
  wire  initBits_7; // @[StoreQueue.scala 70:64:@227.4]
  wire [6:0] _T_1676; // @[util.scala 14:20:@229.4]
  wire [6:0] _T_1677; // @[util.scala 14:20:@230.4]
  wire [5:0] _T_1678; // @[util.scala 14:20:@231.4]
  wire [5:0] _GEN_136; // @[util.scala 14:25:@232.4]
  wire [4:0] _T_1679; // @[util.scala 14:25:@232.4]
  wire  _T_1680; // @[StoreQueue.scala 70:46:@233.4]
  wire  initBits_8; // @[StoreQueue.scala 70:64:@234.4]
  wire [6:0] _T_1685; // @[util.scala 14:20:@236.4]
  wire [6:0] _T_1686; // @[util.scala 14:20:@237.4]
  wire [5:0] _T_1687; // @[util.scala 14:20:@238.4]
  wire [5:0] _GEN_152; // @[util.scala 14:25:@239.4]
  wire [4:0] _T_1688; // @[util.scala 14:25:@239.4]
  wire  _T_1689; // @[StoreQueue.scala 70:46:@240.4]
  wire  initBits_9; // @[StoreQueue.scala 70:64:@241.4]
  wire [6:0] _T_1694; // @[util.scala 14:20:@243.4]
  wire [6:0] _T_1695; // @[util.scala 14:20:@244.4]
  wire [5:0] _T_1696; // @[util.scala 14:20:@245.4]
  wire [5:0] _GEN_170; // @[util.scala 14:25:@246.4]
  wire [4:0] _T_1697; // @[util.scala 14:25:@246.4]
  wire  _T_1698; // @[StoreQueue.scala 70:46:@247.4]
  wire  initBits_10; // @[StoreQueue.scala 70:64:@248.4]
  wire [6:0] _T_1703; // @[util.scala 14:20:@250.4]
  wire [6:0] _T_1704; // @[util.scala 14:20:@251.4]
  wire [5:0] _T_1705; // @[util.scala 14:20:@252.4]
  wire [5:0] _GEN_186; // @[util.scala 14:25:@253.4]
  wire [4:0] _T_1706; // @[util.scala 14:25:@253.4]
  wire  _T_1707; // @[StoreQueue.scala 70:46:@254.4]
  wire  initBits_11; // @[StoreQueue.scala 70:64:@255.4]
  wire [6:0] _T_1712; // @[util.scala 14:20:@257.4]
  wire [6:0] _T_1713; // @[util.scala 14:20:@258.4]
  wire [5:0] _T_1714; // @[util.scala 14:20:@259.4]
  wire [5:0] _GEN_204; // @[util.scala 14:25:@260.4]
  wire [4:0] _T_1715; // @[util.scala 14:25:@260.4]
  wire  _T_1716; // @[StoreQueue.scala 70:46:@261.4]
  wire  initBits_12; // @[StoreQueue.scala 70:64:@262.4]
  wire [6:0] _T_1721; // @[util.scala 14:20:@264.4]
  wire [6:0] _T_1722; // @[util.scala 14:20:@265.4]
  wire [5:0] _T_1723; // @[util.scala 14:20:@266.4]
  wire [5:0] _GEN_220; // @[util.scala 14:25:@267.4]
  wire [4:0] _T_1724; // @[util.scala 14:25:@267.4]
  wire  _T_1725; // @[StoreQueue.scala 70:46:@268.4]
  wire  initBits_13; // @[StoreQueue.scala 70:64:@269.4]
  wire [6:0] _T_1730; // @[util.scala 14:20:@271.4]
  wire [6:0] _T_1731; // @[util.scala 14:20:@272.4]
  wire [5:0] _T_1732; // @[util.scala 14:20:@273.4]
  wire [5:0] _GEN_238; // @[util.scala 14:25:@274.4]
  wire [4:0] _T_1733; // @[util.scala 14:25:@274.4]
  wire  _T_1734; // @[StoreQueue.scala 70:46:@275.4]
  wire  initBits_14; // @[StoreQueue.scala 70:64:@276.4]
  wire [6:0] _T_1739; // @[util.scala 14:20:@278.4]
  wire [6:0] _T_1740; // @[util.scala 14:20:@279.4]
  wire [5:0] _T_1741; // @[util.scala 14:20:@280.4]
  wire [5:0] _GEN_254; // @[util.scala 14:25:@281.4]
  wire [4:0] _T_1742; // @[util.scala 14:25:@281.4]
  wire  _T_1743; // @[StoreQueue.scala 70:46:@282.4]
  wire  initBits_15; // @[StoreQueue.scala 70:64:@283.4]
  wire  _T_1766; // @[StoreQueue.scala 72:78:@301.4]
  wire  _T_1767; // @[StoreQueue.scala 72:78:@302.4]
  wire  _T_1768; // @[StoreQueue.scala 72:78:@303.4]
  wire  _T_1769; // @[StoreQueue.scala 72:78:@304.4]
  wire  _T_1770; // @[StoreQueue.scala 72:78:@305.4]
  wire  _T_1771; // @[StoreQueue.scala 72:78:@306.4]
  wire  _T_1772; // @[StoreQueue.scala 72:78:@307.4]
  wire  _T_1773; // @[StoreQueue.scala 72:78:@308.4]
  wire  _T_1774; // @[StoreQueue.scala 72:78:@309.4]
  wire  _T_1775; // @[StoreQueue.scala 72:78:@310.4]
  wire  _T_1776; // @[StoreQueue.scala 72:78:@311.4]
  wire  _T_1777; // @[StoreQueue.scala 72:78:@312.4]
  wire  _T_1778; // @[StoreQueue.scala 72:78:@313.4]
  wire  _T_1779; // @[StoreQueue.scala 72:78:@314.4]
  wire  _T_1780; // @[StoreQueue.scala 72:78:@315.4]
  wire  _T_1781; // @[StoreQueue.scala 72:78:@316.4]
  wire [3:0] _T_1812; // @[:@356.6]
  wire [3:0] _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_15; // @[StoreQueue.scala 76:20:@357.6]
  wire  _GEN_17; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_18; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_19; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_20; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_21; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_22; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_23; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_24; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_25; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_26; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_27; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_28; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_29; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_30; // @[StoreQueue.scala 77:18:@364.6]
  wire  _GEN_31; // @[StoreQueue.scala 77:18:@364.6]
  wire [3:0] _GEN_32; // @[StoreQueue.scala 75:25:@350.4]
  wire  _GEN_33; // @[StoreQueue.scala 75:25:@350.4]
  wire [3:0] _T_1830; // @[:@372.6]
  wire [3:0] _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_49; // @[StoreQueue.scala 76:20:@373.6]
  wire  _GEN_51; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_52; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_53; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_54; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_55; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_56; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_57; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_58; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_59; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_60; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_61; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_62; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_63; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_64; // @[StoreQueue.scala 77:18:@380.6]
  wire  _GEN_65; // @[StoreQueue.scala 77:18:@380.6]
  wire [3:0] _GEN_66; // @[StoreQueue.scala 75:25:@366.4]
  wire  _GEN_67; // @[StoreQueue.scala 75:25:@366.4]
  wire [3:0] _T_1848; // @[:@388.6]
  wire [3:0] _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_83; // @[StoreQueue.scala 76:20:@389.6]
  wire  _GEN_85; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_86; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_87; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_88; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_89; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_90; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_91; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_92; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_93; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_94; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_95; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_96; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_97; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_98; // @[StoreQueue.scala 77:18:@396.6]
  wire  _GEN_99; // @[StoreQueue.scala 77:18:@396.6]
  wire [3:0] _GEN_100; // @[StoreQueue.scala 75:25:@382.4]
  wire  _GEN_101; // @[StoreQueue.scala 75:25:@382.4]
  wire [3:0] _T_1866; // @[:@404.6]
  wire [3:0] _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_117; // @[StoreQueue.scala 76:20:@405.6]
  wire  _GEN_119; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_120; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_121; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_122; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_123; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_124; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_125; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_126; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_127; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_128; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_129; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_130; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_131; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_132; // @[StoreQueue.scala 77:18:@412.6]
  wire  _GEN_133; // @[StoreQueue.scala 77:18:@412.6]
  wire [3:0] _GEN_134; // @[StoreQueue.scala 75:25:@398.4]
  wire  _GEN_135; // @[StoreQueue.scala 75:25:@398.4]
  wire [3:0] _T_1884; // @[:@420.6]
  wire [3:0] _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_151; // @[StoreQueue.scala 76:20:@421.6]
  wire  _GEN_153; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_154; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_155; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_156; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_157; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_158; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_159; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_160; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_161; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_162; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_163; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_164; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_165; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_166; // @[StoreQueue.scala 77:18:@428.6]
  wire  _GEN_167; // @[StoreQueue.scala 77:18:@428.6]
  wire [3:0] _GEN_168; // @[StoreQueue.scala 75:25:@414.4]
  wire  _GEN_169; // @[StoreQueue.scala 75:25:@414.4]
  wire [3:0] _T_1902; // @[:@436.6]
  wire [3:0] _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_185; // @[StoreQueue.scala 76:20:@437.6]
  wire  _GEN_187; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_188; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_189; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_190; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_191; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_192; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_193; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_194; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_195; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_196; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_197; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_198; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_199; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_200; // @[StoreQueue.scala 77:18:@444.6]
  wire  _GEN_201; // @[StoreQueue.scala 77:18:@444.6]
  wire [3:0] _GEN_202; // @[StoreQueue.scala 75:25:@430.4]
  wire  _GEN_203; // @[StoreQueue.scala 75:25:@430.4]
  wire [3:0] _T_1920; // @[:@452.6]
  wire [3:0] _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_219; // @[StoreQueue.scala 76:20:@453.6]
  wire  _GEN_221; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_222; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_223; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_224; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_225; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_226; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_227; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_228; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_229; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_230; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_231; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_232; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_233; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_234; // @[StoreQueue.scala 77:18:@460.6]
  wire  _GEN_235; // @[StoreQueue.scala 77:18:@460.6]
  wire [3:0] _GEN_236; // @[StoreQueue.scala 75:25:@446.4]
  wire  _GEN_237; // @[StoreQueue.scala 75:25:@446.4]
  wire [3:0] _T_1938; // @[:@468.6]
  wire [3:0] _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_253; // @[StoreQueue.scala 76:20:@469.6]
  wire  _GEN_255; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_256; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_257; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_258; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_259; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_260; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_261; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_262; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_263; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_264; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_265; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_266; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_267; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_268; // @[StoreQueue.scala 77:18:@476.6]
  wire  _GEN_269; // @[StoreQueue.scala 77:18:@476.6]
  wire [3:0] _GEN_270; // @[StoreQueue.scala 75:25:@462.4]
  wire  _GEN_271; // @[StoreQueue.scala 75:25:@462.4]
  wire [3:0] _T_1956; // @[:@484.6]
  wire [3:0] _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_287; // @[StoreQueue.scala 76:20:@485.6]
  wire  _GEN_289; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_290; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_291; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_292; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_293; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_294; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_295; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_296; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_297; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_298; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_299; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_300; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_301; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_302; // @[StoreQueue.scala 77:18:@492.6]
  wire  _GEN_303; // @[StoreQueue.scala 77:18:@492.6]
  wire [3:0] _GEN_304; // @[StoreQueue.scala 75:25:@478.4]
  wire  _GEN_305; // @[StoreQueue.scala 75:25:@478.4]
  wire [3:0] _T_1974; // @[:@500.6]
  wire [3:0] _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_321; // @[StoreQueue.scala 76:20:@501.6]
  wire  _GEN_323; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_324; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_325; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_326; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_327; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_328; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_329; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_330; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_331; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_332; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_333; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_334; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_335; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_336; // @[StoreQueue.scala 77:18:@508.6]
  wire  _GEN_337; // @[StoreQueue.scala 77:18:@508.6]
  wire [3:0] _GEN_338; // @[StoreQueue.scala 75:25:@494.4]
  wire  _GEN_339; // @[StoreQueue.scala 75:25:@494.4]
  wire [3:0] _T_1992; // @[:@516.6]
  wire [3:0] _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_355; // @[StoreQueue.scala 76:20:@517.6]
  wire  _GEN_357; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_358; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_359; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_360; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_361; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_362; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_363; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_364; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_365; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_366; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_367; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_368; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_369; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_370; // @[StoreQueue.scala 77:18:@524.6]
  wire  _GEN_371; // @[StoreQueue.scala 77:18:@524.6]
  wire [3:0] _GEN_372; // @[StoreQueue.scala 75:25:@510.4]
  wire  _GEN_373; // @[StoreQueue.scala 75:25:@510.4]
  wire [3:0] _T_2010; // @[:@532.6]
  wire [3:0] _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_389; // @[StoreQueue.scala 76:20:@533.6]
  wire  _GEN_391; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_392; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_393; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_394; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_395; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_396; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_397; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_398; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_399; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_400; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_401; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_402; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_403; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_404; // @[StoreQueue.scala 77:18:@540.6]
  wire  _GEN_405; // @[StoreQueue.scala 77:18:@540.6]
  wire [3:0] _GEN_406; // @[StoreQueue.scala 75:25:@526.4]
  wire  _GEN_407; // @[StoreQueue.scala 75:25:@526.4]
  wire [3:0] _T_2028; // @[:@548.6]
  wire [3:0] _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_423; // @[StoreQueue.scala 76:20:@549.6]
  wire  _GEN_425; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_426; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_427; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_428; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_429; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_430; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_431; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_432; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_433; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_434; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_435; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_436; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_437; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_438; // @[StoreQueue.scala 77:18:@556.6]
  wire  _GEN_439; // @[StoreQueue.scala 77:18:@556.6]
  wire [3:0] _GEN_440; // @[StoreQueue.scala 75:25:@542.4]
  wire  _GEN_441; // @[StoreQueue.scala 75:25:@542.4]
  wire [3:0] _T_2046; // @[:@564.6]
  wire [3:0] _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_457; // @[StoreQueue.scala 76:20:@565.6]
  wire  _GEN_459; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_460; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_461; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_462; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_463; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_464; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_465; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_466; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_467; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_468; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_469; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_470; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_471; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_472; // @[StoreQueue.scala 77:18:@572.6]
  wire  _GEN_473; // @[StoreQueue.scala 77:18:@572.6]
  wire [3:0] _GEN_474; // @[StoreQueue.scala 75:25:@558.4]
  wire  _GEN_475; // @[StoreQueue.scala 75:25:@558.4]
  wire [3:0] _T_2064; // @[:@580.6]
  wire [3:0] _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_491; // @[StoreQueue.scala 76:20:@581.6]
  wire  _GEN_493; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_494; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_495; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_496; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_497; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_498; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_499; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_500; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_501; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_502; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_503; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_504; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_505; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_506; // @[StoreQueue.scala 77:18:@588.6]
  wire  _GEN_507; // @[StoreQueue.scala 77:18:@588.6]
  wire [3:0] _GEN_508; // @[StoreQueue.scala 75:25:@574.4]
  wire  _GEN_509; // @[StoreQueue.scala 75:25:@574.4]
  wire [3:0] _T_2082; // @[:@596.6]
  wire [3:0] _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_525; // @[StoreQueue.scala 76:20:@597.6]
  wire  _GEN_527; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_528; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_529; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_530; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_531; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_532; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_533; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_534; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_535; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_536; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_537; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_538; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_539; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_540; // @[StoreQueue.scala 77:18:@604.6]
  wire  _GEN_541; // @[StoreQueue.scala 77:18:@604.6]
  wire [3:0] _GEN_542; // @[StoreQueue.scala 75:25:@590.4]
  wire  _GEN_543; // @[StoreQueue.scala 75:25:@590.4]
  reg [3:0] previousLoadHead; // @[StoreQueue.scala 92:33:@606.4]
  reg [31:0] _RAND_146;
  wire [4:0] _T_2104; // @[util.scala 10:8:@615.6]
  wire [4:0] _GEN_272; // @[util.scala 10:14:@616.6]
  wire [4:0] _T_2105; // @[util.scala 10:14:@616.6]
  wire [4:0] _GEN_1267; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2106; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2107; // @[StoreQueue.scala 95:50:@618.6]
  wire  _T_2109; // @[StoreQueue.scala 95:35:@619.6]
  wire  _T_2111; // @[StoreQueue.scala 100:35:@627.8]
  wire  _T_2112; // @[StoreQueue.scala 100:87:@628.8]
  wire  _T_2113; // @[StoreQueue.scala 100:61:@629.8]
  wire  _T_2115; // @[StoreQueue.scala 102:35:@634.10]
  wire  _T_2116; // @[StoreQueue.scala 103:23:@635.10]
  wire  _T_2117; // @[StoreQueue.scala 103:75:@636.10]
  wire  _T_2118; // @[StoreQueue.scala 103:49:@637.10]
  wire  _T_2120; // @[StoreQueue.scala 103:9:@638.10]
  wire  _T_2121; // @[StoreQueue.scala 102:49:@639.10]
  wire  _GEN_560; // @[StoreQueue.scala 103:96:@640.10]
  wire  _GEN_561; // @[StoreQueue.scala 100:102:@630.8]
  wire  _GEN_562; // @[StoreQueue.scala 98:26:@623.6]
  wire  _GEN_563; // @[StoreQueue.scala 94:35:@608.4]
  wire [4:0] _T_2134; // @[util.scala 10:8:@651.6]
  wire [4:0] _GEN_288; // @[util.scala 10:14:@652.6]
  wire [4:0] _T_2135; // @[util.scala 10:14:@652.6]
  wire  _T_2136; // @[StoreQueue.scala 96:56:@653.6]
  wire  _T_2137; // @[StoreQueue.scala 95:50:@654.6]
  wire  _T_2139; // @[StoreQueue.scala 95:35:@655.6]
  wire  _T_2141; // @[StoreQueue.scala 100:35:@663.8]
  wire  _T_2142; // @[StoreQueue.scala 100:87:@664.8]
  wire  _T_2143; // @[StoreQueue.scala 100:61:@665.8]
  wire  _T_2146; // @[StoreQueue.scala 103:23:@671.10]
  wire  _T_2147; // @[StoreQueue.scala 103:75:@672.10]
  wire  _T_2148; // @[StoreQueue.scala 103:49:@673.10]
  wire  _T_2150; // @[StoreQueue.scala 103:9:@674.10]
  wire  _T_2151; // @[StoreQueue.scala 102:49:@675.10]
  wire  _GEN_580; // @[StoreQueue.scala 103:96:@676.10]
  wire  _GEN_581; // @[StoreQueue.scala 100:102:@666.8]
  wire  _GEN_582; // @[StoreQueue.scala 98:26:@659.6]
  wire  _GEN_583; // @[StoreQueue.scala 94:35:@644.4]
  wire [4:0] _T_2164; // @[util.scala 10:8:@687.6]
  wire [4:0] _GEN_306; // @[util.scala 10:14:@688.6]
  wire [4:0] _T_2165; // @[util.scala 10:14:@688.6]
  wire  _T_2166; // @[StoreQueue.scala 96:56:@689.6]
  wire  _T_2167; // @[StoreQueue.scala 95:50:@690.6]
  wire  _T_2169; // @[StoreQueue.scala 95:35:@691.6]
  wire  _T_2171; // @[StoreQueue.scala 100:35:@699.8]
  wire  _T_2172; // @[StoreQueue.scala 100:87:@700.8]
  wire  _T_2173; // @[StoreQueue.scala 100:61:@701.8]
  wire  _T_2176; // @[StoreQueue.scala 103:23:@707.10]
  wire  _T_2177; // @[StoreQueue.scala 103:75:@708.10]
  wire  _T_2178; // @[StoreQueue.scala 103:49:@709.10]
  wire  _T_2180; // @[StoreQueue.scala 103:9:@710.10]
  wire  _T_2181; // @[StoreQueue.scala 102:49:@711.10]
  wire  _GEN_600; // @[StoreQueue.scala 103:96:@712.10]
  wire  _GEN_601; // @[StoreQueue.scala 100:102:@702.8]
  wire  _GEN_602; // @[StoreQueue.scala 98:26:@695.6]
  wire  _GEN_603; // @[StoreQueue.scala 94:35:@680.4]
  wire [4:0] _T_2194; // @[util.scala 10:8:@723.6]
  wire [4:0] _GEN_322; // @[util.scala 10:14:@724.6]
  wire [4:0] _T_2195; // @[util.scala 10:14:@724.6]
  wire  _T_2196; // @[StoreQueue.scala 96:56:@725.6]
  wire  _T_2197; // @[StoreQueue.scala 95:50:@726.6]
  wire  _T_2199; // @[StoreQueue.scala 95:35:@727.6]
  wire  _T_2201; // @[StoreQueue.scala 100:35:@735.8]
  wire  _T_2202; // @[StoreQueue.scala 100:87:@736.8]
  wire  _T_2203; // @[StoreQueue.scala 100:61:@737.8]
  wire  _T_2206; // @[StoreQueue.scala 103:23:@743.10]
  wire  _T_2207; // @[StoreQueue.scala 103:75:@744.10]
  wire  _T_2208; // @[StoreQueue.scala 103:49:@745.10]
  wire  _T_2210; // @[StoreQueue.scala 103:9:@746.10]
  wire  _T_2211; // @[StoreQueue.scala 102:49:@747.10]
  wire  _GEN_620; // @[StoreQueue.scala 103:96:@748.10]
  wire  _GEN_621; // @[StoreQueue.scala 100:102:@738.8]
  wire  _GEN_622; // @[StoreQueue.scala 98:26:@731.6]
  wire  _GEN_623; // @[StoreQueue.scala 94:35:@716.4]
  wire [4:0] _T_2224; // @[util.scala 10:8:@759.6]
  wire [4:0] _GEN_340; // @[util.scala 10:14:@760.6]
  wire [4:0] _T_2225; // @[util.scala 10:14:@760.6]
  wire  _T_2226; // @[StoreQueue.scala 96:56:@761.6]
  wire  _T_2227; // @[StoreQueue.scala 95:50:@762.6]
  wire  _T_2229; // @[StoreQueue.scala 95:35:@763.6]
  wire  _T_2231; // @[StoreQueue.scala 100:35:@771.8]
  wire  _T_2232; // @[StoreQueue.scala 100:87:@772.8]
  wire  _T_2233; // @[StoreQueue.scala 100:61:@773.8]
  wire  _T_2236; // @[StoreQueue.scala 103:23:@779.10]
  wire  _T_2237; // @[StoreQueue.scala 103:75:@780.10]
  wire  _T_2238; // @[StoreQueue.scala 103:49:@781.10]
  wire  _T_2240; // @[StoreQueue.scala 103:9:@782.10]
  wire  _T_2241; // @[StoreQueue.scala 102:49:@783.10]
  wire  _GEN_640; // @[StoreQueue.scala 103:96:@784.10]
  wire  _GEN_641; // @[StoreQueue.scala 100:102:@774.8]
  wire  _GEN_642; // @[StoreQueue.scala 98:26:@767.6]
  wire  _GEN_643; // @[StoreQueue.scala 94:35:@752.4]
  wire [4:0] _T_2254; // @[util.scala 10:8:@795.6]
  wire [4:0] _GEN_356; // @[util.scala 10:14:@796.6]
  wire [4:0] _T_2255; // @[util.scala 10:14:@796.6]
  wire  _T_2256; // @[StoreQueue.scala 96:56:@797.6]
  wire  _T_2257; // @[StoreQueue.scala 95:50:@798.6]
  wire  _T_2259; // @[StoreQueue.scala 95:35:@799.6]
  wire  _T_2261; // @[StoreQueue.scala 100:35:@807.8]
  wire  _T_2262; // @[StoreQueue.scala 100:87:@808.8]
  wire  _T_2263; // @[StoreQueue.scala 100:61:@809.8]
  wire  _T_2266; // @[StoreQueue.scala 103:23:@815.10]
  wire  _T_2267; // @[StoreQueue.scala 103:75:@816.10]
  wire  _T_2268; // @[StoreQueue.scala 103:49:@817.10]
  wire  _T_2270; // @[StoreQueue.scala 103:9:@818.10]
  wire  _T_2271; // @[StoreQueue.scala 102:49:@819.10]
  wire  _GEN_660; // @[StoreQueue.scala 103:96:@820.10]
  wire  _GEN_661; // @[StoreQueue.scala 100:102:@810.8]
  wire  _GEN_662; // @[StoreQueue.scala 98:26:@803.6]
  wire  _GEN_663; // @[StoreQueue.scala 94:35:@788.4]
  wire [4:0] _T_2284; // @[util.scala 10:8:@831.6]
  wire [4:0] _GEN_374; // @[util.scala 10:14:@832.6]
  wire [4:0] _T_2285; // @[util.scala 10:14:@832.6]
  wire  _T_2286; // @[StoreQueue.scala 96:56:@833.6]
  wire  _T_2287; // @[StoreQueue.scala 95:50:@834.6]
  wire  _T_2289; // @[StoreQueue.scala 95:35:@835.6]
  wire  _T_2291; // @[StoreQueue.scala 100:35:@843.8]
  wire  _T_2292; // @[StoreQueue.scala 100:87:@844.8]
  wire  _T_2293; // @[StoreQueue.scala 100:61:@845.8]
  wire  _T_2296; // @[StoreQueue.scala 103:23:@851.10]
  wire  _T_2297; // @[StoreQueue.scala 103:75:@852.10]
  wire  _T_2298; // @[StoreQueue.scala 103:49:@853.10]
  wire  _T_2300; // @[StoreQueue.scala 103:9:@854.10]
  wire  _T_2301; // @[StoreQueue.scala 102:49:@855.10]
  wire  _GEN_680; // @[StoreQueue.scala 103:96:@856.10]
  wire  _GEN_681; // @[StoreQueue.scala 100:102:@846.8]
  wire  _GEN_682; // @[StoreQueue.scala 98:26:@839.6]
  wire  _GEN_683; // @[StoreQueue.scala 94:35:@824.4]
  wire [4:0] _T_2314; // @[util.scala 10:8:@867.6]
  wire [4:0] _GEN_390; // @[util.scala 10:14:@868.6]
  wire [4:0] _T_2315; // @[util.scala 10:14:@868.6]
  wire  _T_2316; // @[StoreQueue.scala 96:56:@869.6]
  wire  _T_2317; // @[StoreQueue.scala 95:50:@870.6]
  wire  _T_2319; // @[StoreQueue.scala 95:35:@871.6]
  wire  _T_2321; // @[StoreQueue.scala 100:35:@879.8]
  wire  _T_2322; // @[StoreQueue.scala 100:87:@880.8]
  wire  _T_2323; // @[StoreQueue.scala 100:61:@881.8]
  wire  _T_2326; // @[StoreQueue.scala 103:23:@887.10]
  wire  _T_2327; // @[StoreQueue.scala 103:75:@888.10]
  wire  _T_2328; // @[StoreQueue.scala 103:49:@889.10]
  wire  _T_2330; // @[StoreQueue.scala 103:9:@890.10]
  wire  _T_2331; // @[StoreQueue.scala 102:49:@891.10]
  wire  _GEN_700; // @[StoreQueue.scala 103:96:@892.10]
  wire  _GEN_701; // @[StoreQueue.scala 100:102:@882.8]
  wire  _GEN_702; // @[StoreQueue.scala 98:26:@875.6]
  wire  _GEN_703; // @[StoreQueue.scala 94:35:@860.4]
  wire [4:0] _T_2344; // @[util.scala 10:8:@903.6]
  wire [4:0] _GEN_408; // @[util.scala 10:14:@904.6]
  wire [4:0] _T_2345; // @[util.scala 10:14:@904.6]
  wire  _T_2346; // @[StoreQueue.scala 96:56:@905.6]
  wire  _T_2347; // @[StoreQueue.scala 95:50:@906.6]
  wire  _T_2349; // @[StoreQueue.scala 95:35:@907.6]
  wire  _T_2351; // @[StoreQueue.scala 100:35:@915.8]
  wire  _T_2352; // @[StoreQueue.scala 100:87:@916.8]
  wire  _T_2353; // @[StoreQueue.scala 100:61:@917.8]
  wire  _T_2356; // @[StoreQueue.scala 103:23:@923.10]
  wire  _T_2357; // @[StoreQueue.scala 103:75:@924.10]
  wire  _T_2358; // @[StoreQueue.scala 103:49:@925.10]
  wire  _T_2360; // @[StoreQueue.scala 103:9:@926.10]
  wire  _T_2361; // @[StoreQueue.scala 102:49:@927.10]
  wire  _GEN_720; // @[StoreQueue.scala 103:96:@928.10]
  wire  _GEN_721; // @[StoreQueue.scala 100:102:@918.8]
  wire  _GEN_722; // @[StoreQueue.scala 98:26:@911.6]
  wire  _GEN_723; // @[StoreQueue.scala 94:35:@896.4]
  wire [4:0] _T_2374; // @[util.scala 10:8:@939.6]
  wire [4:0] _GEN_424; // @[util.scala 10:14:@940.6]
  wire [4:0] _T_2375; // @[util.scala 10:14:@940.6]
  wire  _T_2376; // @[StoreQueue.scala 96:56:@941.6]
  wire  _T_2377; // @[StoreQueue.scala 95:50:@942.6]
  wire  _T_2379; // @[StoreQueue.scala 95:35:@943.6]
  wire  _T_2381; // @[StoreQueue.scala 100:35:@951.8]
  wire  _T_2382; // @[StoreQueue.scala 100:87:@952.8]
  wire  _T_2383; // @[StoreQueue.scala 100:61:@953.8]
  wire  _T_2386; // @[StoreQueue.scala 103:23:@959.10]
  wire  _T_2387; // @[StoreQueue.scala 103:75:@960.10]
  wire  _T_2388; // @[StoreQueue.scala 103:49:@961.10]
  wire  _T_2390; // @[StoreQueue.scala 103:9:@962.10]
  wire  _T_2391; // @[StoreQueue.scala 102:49:@963.10]
  wire  _GEN_740; // @[StoreQueue.scala 103:96:@964.10]
  wire  _GEN_741; // @[StoreQueue.scala 100:102:@954.8]
  wire  _GEN_742; // @[StoreQueue.scala 98:26:@947.6]
  wire  _GEN_743; // @[StoreQueue.scala 94:35:@932.4]
  wire [4:0] _T_2404; // @[util.scala 10:8:@975.6]
  wire [4:0] _GEN_442; // @[util.scala 10:14:@976.6]
  wire [4:0] _T_2405; // @[util.scala 10:14:@976.6]
  wire  _T_2406; // @[StoreQueue.scala 96:56:@977.6]
  wire  _T_2407; // @[StoreQueue.scala 95:50:@978.6]
  wire  _T_2409; // @[StoreQueue.scala 95:35:@979.6]
  wire  _T_2411; // @[StoreQueue.scala 100:35:@987.8]
  wire  _T_2412; // @[StoreQueue.scala 100:87:@988.8]
  wire  _T_2413; // @[StoreQueue.scala 100:61:@989.8]
  wire  _T_2416; // @[StoreQueue.scala 103:23:@995.10]
  wire  _T_2417; // @[StoreQueue.scala 103:75:@996.10]
  wire  _T_2418; // @[StoreQueue.scala 103:49:@997.10]
  wire  _T_2420; // @[StoreQueue.scala 103:9:@998.10]
  wire  _T_2421; // @[StoreQueue.scala 102:49:@999.10]
  wire  _GEN_760; // @[StoreQueue.scala 103:96:@1000.10]
  wire  _GEN_761; // @[StoreQueue.scala 100:102:@990.8]
  wire  _GEN_762; // @[StoreQueue.scala 98:26:@983.6]
  wire  _GEN_763; // @[StoreQueue.scala 94:35:@968.4]
  wire [4:0] _T_2434; // @[util.scala 10:8:@1011.6]
  wire [4:0] _GEN_458; // @[util.scala 10:14:@1012.6]
  wire [4:0] _T_2435; // @[util.scala 10:14:@1012.6]
  wire  _T_2436; // @[StoreQueue.scala 96:56:@1013.6]
  wire  _T_2437; // @[StoreQueue.scala 95:50:@1014.6]
  wire  _T_2439; // @[StoreQueue.scala 95:35:@1015.6]
  wire  _T_2441; // @[StoreQueue.scala 100:35:@1023.8]
  wire  _T_2442; // @[StoreQueue.scala 100:87:@1024.8]
  wire  _T_2443; // @[StoreQueue.scala 100:61:@1025.8]
  wire  _T_2446; // @[StoreQueue.scala 103:23:@1031.10]
  wire  _T_2447; // @[StoreQueue.scala 103:75:@1032.10]
  wire  _T_2448; // @[StoreQueue.scala 103:49:@1033.10]
  wire  _T_2450; // @[StoreQueue.scala 103:9:@1034.10]
  wire  _T_2451; // @[StoreQueue.scala 102:49:@1035.10]
  wire  _GEN_780; // @[StoreQueue.scala 103:96:@1036.10]
  wire  _GEN_781; // @[StoreQueue.scala 100:102:@1026.8]
  wire  _GEN_782; // @[StoreQueue.scala 98:26:@1019.6]
  wire  _GEN_783; // @[StoreQueue.scala 94:35:@1004.4]
  wire [4:0] _T_2464; // @[util.scala 10:8:@1047.6]
  wire [4:0] _GEN_476; // @[util.scala 10:14:@1048.6]
  wire [4:0] _T_2465; // @[util.scala 10:14:@1048.6]
  wire  _T_2466; // @[StoreQueue.scala 96:56:@1049.6]
  wire  _T_2467; // @[StoreQueue.scala 95:50:@1050.6]
  wire  _T_2469; // @[StoreQueue.scala 95:35:@1051.6]
  wire  _T_2471; // @[StoreQueue.scala 100:35:@1059.8]
  wire  _T_2472; // @[StoreQueue.scala 100:87:@1060.8]
  wire  _T_2473; // @[StoreQueue.scala 100:61:@1061.8]
  wire  _T_2476; // @[StoreQueue.scala 103:23:@1067.10]
  wire  _T_2477; // @[StoreQueue.scala 103:75:@1068.10]
  wire  _T_2478; // @[StoreQueue.scala 103:49:@1069.10]
  wire  _T_2480; // @[StoreQueue.scala 103:9:@1070.10]
  wire  _T_2481; // @[StoreQueue.scala 102:49:@1071.10]
  wire  _GEN_800; // @[StoreQueue.scala 103:96:@1072.10]
  wire  _GEN_801; // @[StoreQueue.scala 100:102:@1062.8]
  wire  _GEN_802; // @[StoreQueue.scala 98:26:@1055.6]
  wire  _GEN_803; // @[StoreQueue.scala 94:35:@1040.4]
  wire [4:0] _T_2494; // @[util.scala 10:8:@1083.6]
  wire [4:0] _GEN_492; // @[util.scala 10:14:@1084.6]
  wire [4:0] _T_2495; // @[util.scala 10:14:@1084.6]
  wire  _T_2496; // @[StoreQueue.scala 96:56:@1085.6]
  wire  _T_2497; // @[StoreQueue.scala 95:50:@1086.6]
  wire  _T_2499; // @[StoreQueue.scala 95:35:@1087.6]
  wire  _T_2501; // @[StoreQueue.scala 100:35:@1095.8]
  wire  _T_2502; // @[StoreQueue.scala 100:87:@1096.8]
  wire  _T_2503; // @[StoreQueue.scala 100:61:@1097.8]
  wire  _T_2506; // @[StoreQueue.scala 103:23:@1103.10]
  wire  _T_2507; // @[StoreQueue.scala 103:75:@1104.10]
  wire  _T_2508; // @[StoreQueue.scala 103:49:@1105.10]
  wire  _T_2510; // @[StoreQueue.scala 103:9:@1106.10]
  wire  _T_2511; // @[StoreQueue.scala 102:49:@1107.10]
  wire  _GEN_820; // @[StoreQueue.scala 103:96:@1108.10]
  wire  _GEN_821; // @[StoreQueue.scala 100:102:@1098.8]
  wire  _GEN_822; // @[StoreQueue.scala 98:26:@1091.6]
  wire  _GEN_823; // @[StoreQueue.scala 94:35:@1076.4]
  wire [4:0] _T_2524; // @[util.scala 10:8:@1119.6]
  wire [4:0] _GEN_510; // @[util.scala 10:14:@1120.6]
  wire [4:0] _T_2525; // @[util.scala 10:14:@1120.6]
  wire  _T_2526; // @[StoreQueue.scala 96:56:@1121.6]
  wire  _T_2527; // @[StoreQueue.scala 95:50:@1122.6]
  wire  _T_2529; // @[StoreQueue.scala 95:35:@1123.6]
  wire  _T_2531; // @[StoreQueue.scala 100:35:@1131.8]
  wire  _T_2532; // @[StoreQueue.scala 100:87:@1132.8]
  wire  _T_2533; // @[StoreQueue.scala 100:61:@1133.8]
  wire  _T_2536; // @[StoreQueue.scala 103:23:@1139.10]
  wire  _T_2537; // @[StoreQueue.scala 103:75:@1140.10]
  wire  _T_2538; // @[StoreQueue.scala 103:49:@1141.10]
  wire  _T_2540; // @[StoreQueue.scala 103:9:@1142.10]
  wire  _T_2541; // @[StoreQueue.scala 102:49:@1143.10]
  wire  _GEN_840; // @[StoreQueue.scala 103:96:@1144.10]
  wire  _GEN_841; // @[StoreQueue.scala 100:102:@1134.8]
  wire  _GEN_842; // @[StoreQueue.scala 98:26:@1127.6]
  wire  _GEN_843; // @[StoreQueue.scala 94:35:@1112.4]
  wire [4:0] _T_2554; // @[util.scala 10:8:@1155.6]
  wire [4:0] _GEN_526; // @[util.scala 10:14:@1156.6]
  wire [4:0] _T_2555; // @[util.scala 10:14:@1156.6]
  wire  _T_2556; // @[StoreQueue.scala 96:56:@1157.6]
  wire  _T_2557; // @[StoreQueue.scala 95:50:@1158.6]
  wire  _T_2559; // @[StoreQueue.scala 95:35:@1159.6]
  wire  _T_2561; // @[StoreQueue.scala 100:35:@1167.8]
  wire  _T_2562; // @[StoreQueue.scala 100:87:@1168.8]
  wire  _T_2563; // @[StoreQueue.scala 100:61:@1169.8]
  wire  _T_2566; // @[StoreQueue.scala 103:23:@1175.10]
  wire  _T_2567; // @[StoreQueue.scala 103:75:@1176.10]
  wire  _T_2568; // @[StoreQueue.scala 103:49:@1177.10]
  wire  _T_2570; // @[StoreQueue.scala 103:9:@1178.10]
  wire  _T_2571; // @[StoreQueue.scala 102:49:@1179.10]
  wire  _GEN_860; // @[StoreQueue.scala 103:96:@1180.10]
  wire  _GEN_861; // @[StoreQueue.scala 100:102:@1170.8]
  wire  _GEN_862; // @[StoreQueue.scala 98:26:@1163.6]
  wire  _GEN_863; // @[StoreQueue.scala 94:35:@1148.4]
  wire  _T_2573; // @[StoreQueue.scala 119:103:@1184.4]
  wire  _T_2575; // @[StoreQueue.scala 120:17:@1185.4]
  wire  _T_2577; // @[StoreQueue.scala 120:35:@1186.4]
  wire  _T_2578; // @[StoreQueue.scala 120:26:@1187.4]
  wire  _T_2580; // @[StoreQueue.scala 120:50:@1188.4]
  wire  _T_2582; // @[StoreQueue.scala 120:81:@1189.4]
  wire  _T_2584; // @[StoreQueue.scala 120:99:@1190.4]
  wire  _T_2585; // @[StoreQueue.scala 120:90:@1191.4]
  wire  _T_2587; // @[StoreQueue.scala 120:67:@1192.4]
  wire  _T_2588; // @[StoreQueue.scala 120:64:@1193.4]
  wire  validEntriesInLoadQ_0; // @[StoreQueue.scala 119:90:@1194.4]
  wire  _T_2592; // @[StoreQueue.scala 120:17:@1196.4]
  wire  _T_2594; // @[StoreQueue.scala 120:35:@1197.4]
  wire  _T_2595; // @[StoreQueue.scala 120:26:@1198.4]
  wire  _T_2599; // @[StoreQueue.scala 120:81:@1200.4]
  wire  _T_2601; // @[StoreQueue.scala 120:99:@1201.4]
  wire  _T_2602; // @[StoreQueue.scala 120:90:@1202.4]
  wire  _T_2604; // @[StoreQueue.scala 120:67:@1203.4]
  wire  _T_2605; // @[StoreQueue.scala 120:64:@1204.4]
  wire  validEntriesInLoadQ_1; // @[StoreQueue.scala 119:90:@1205.4]
  wire  _T_2609; // @[StoreQueue.scala 120:17:@1207.4]
  wire  _T_2611; // @[StoreQueue.scala 120:35:@1208.4]
  wire  _T_2612; // @[StoreQueue.scala 120:26:@1209.4]
  wire  _T_2616; // @[StoreQueue.scala 120:81:@1211.4]
  wire  _T_2618; // @[StoreQueue.scala 120:99:@1212.4]
  wire  _T_2619; // @[StoreQueue.scala 120:90:@1213.4]
  wire  _T_2621; // @[StoreQueue.scala 120:67:@1214.4]
  wire  _T_2622; // @[StoreQueue.scala 120:64:@1215.4]
  wire  validEntriesInLoadQ_2; // @[StoreQueue.scala 119:90:@1216.4]
  wire  _T_2626; // @[StoreQueue.scala 120:17:@1218.4]
  wire  _T_2628; // @[StoreQueue.scala 120:35:@1219.4]
  wire  _T_2629; // @[StoreQueue.scala 120:26:@1220.4]
  wire  _T_2633; // @[StoreQueue.scala 120:81:@1222.4]
  wire  _T_2635; // @[StoreQueue.scala 120:99:@1223.4]
  wire  _T_2636; // @[StoreQueue.scala 120:90:@1224.4]
  wire  _T_2638; // @[StoreQueue.scala 120:67:@1225.4]
  wire  _T_2639; // @[StoreQueue.scala 120:64:@1226.4]
  wire  validEntriesInLoadQ_3; // @[StoreQueue.scala 119:90:@1227.4]
  wire  _T_2643; // @[StoreQueue.scala 120:17:@1229.4]
  wire  _T_2645; // @[StoreQueue.scala 120:35:@1230.4]
  wire  _T_2646; // @[StoreQueue.scala 120:26:@1231.4]
  wire  _T_2650; // @[StoreQueue.scala 120:81:@1233.4]
  wire  _T_2652; // @[StoreQueue.scala 120:99:@1234.4]
  wire  _T_2653; // @[StoreQueue.scala 120:90:@1235.4]
  wire  _T_2655; // @[StoreQueue.scala 120:67:@1236.4]
  wire  _T_2656; // @[StoreQueue.scala 120:64:@1237.4]
  wire  validEntriesInLoadQ_4; // @[StoreQueue.scala 119:90:@1238.4]
  wire  _T_2660; // @[StoreQueue.scala 120:17:@1240.4]
  wire  _T_2662; // @[StoreQueue.scala 120:35:@1241.4]
  wire  _T_2663; // @[StoreQueue.scala 120:26:@1242.4]
  wire  _T_2667; // @[StoreQueue.scala 120:81:@1244.4]
  wire  _T_2669; // @[StoreQueue.scala 120:99:@1245.4]
  wire  _T_2670; // @[StoreQueue.scala 120:90:@1246.4]
  wire  _T_2672; // @[StoreQueue.scala 120:67:@1247.4]
  wire  _T_2673; // @[StoreQueue.scala 120:64:@1248.4]
  wire  validEntriesInLoadQ_5; // @[StoreQueue.scala 119:90:@1249.4]
  wire  _T_2677; // @[StoreQueue.scala 120:17:@1251.4]
  wire  _T_2679; // @[StoreQueue.scala 120:35:@1252.4]
  wire  _T_2680; // @[StoreQueue.scala 120:26:@1253.4]
  wire  _T_2684; // @[StoreQueue.scala 120:81:@1255.4]
  wire  _T_2686; // @[StoreQueue.scala 120:99:@1256.4]
  wire  _T_2687; // @[StoreQueue.scala 120:90:@1257.4]
  wire  _T_2689; // @[StoreQueue.scala 120:67:@1258.4]
  wire  _T_2690; // @[StoreQueue.scala 120:64:@1259.4]
  wire  validEntriesInLoadQ_6; // @[StoreQueue.scala 119:90:@1260.4]
  wire  _T_2694; // @[StoreQueue.scala 120:17:@1262.4]
  wire  _T_2696; // @[StoreQueue.scala 120:35:@1263.4]
  wire  _T_2697; // @[StoreQueue.scala 120:26:@1264.4]
  wire  _T_2701; // @[StoreQueue.scala 120:81:@1266.4]
  wire  _T_2703; // @[StoreQueue.scala 120:99:@1267.4]
  wire  _T_2704; // @[StoreQueue.scala 120:90:@1268.4]
  wire  _T_2706; // @[StoreQueue.scala 120:67:@1269.4]
  wire  _T_2707; // @[StoreQueue.scala 120:64:@1270.4]
  wire  validEntriesInLoadQ_7; // @[StoreQueue.scala 119:90:@1271.4]
  wire  _T_2711; // @[StoreQueue.scala 120:17:@1273.4]
  wire  _T_2713; // @[StoreQueue.scala 120:35:@1274.4]
  wire  _T_2714; // @[StoreQueue.scala 120:26:@1275.4]
  wire  _T_2718; // @[StoreQueue.scala 120:81:@1277.4]
  wire  _T_2720; // @[StoreQueue.scala 120:99:@1278.4]
  wire  _T_2721; // @[StoreQueue.scala 120:90:@1279.4]
  wire  _T_2723; // @[StoreQueue.scala 120:67:@1280.4]
  wire  _T_2724; // @[StoreQueue.scala 120:64:@1281.4]
  wire  validEntriesInLoadQ_8; // @[StoreQueue.scala 119:90:@1282.4]
  wire  _T_2728; // @[StoreQueue.scala 120:17:@1284.4]
  wire  _T_2730; // @[StoreQueue.scala 120:35:@1285.4]
  wire  _T_2731; // @[StoreQueue.scala 120:26:@1286.4]
  wire  _T_2735; // @[StoreQueue.scala 120:81:@1288.4]
  wire  _T_2737; // @[StoreQueue.scala 120:99:@1289.4]
  wire  _T_2738; // @[StoreQueue.scala 120:90:@1290.4]
  wire  _T_2740; // @[StoreQueue.scala 120:67:@1291.4]
  wire  _T_2741; // @[StoreQueue.scala 120:64:@1292.4]
  wire  validEntriesInLoadQ_9; // @[StoreQueue.scala 119:90:@1293.4]
  wire  _T_2745; // @[StoreQueue.scala 120:17:@1295.4]
  wire  _T_2747; // @[StoreQueue.scala 120:35:@1296.4]
  wire  _T_2748; // @[StoreQueue.scala 120:26:@1297.4]
  wire  _T_2752; // @[StoreQueue.scala 120:81:@1299.4]
  wire  _T_2754; // @[StoreQueue.scala 120:99:@1300.4]
  wire  _T_2755; // @[StoreQueue.scala 120:90:@1301.4]
  wire  _T_2757; // @[StoreQueue.scala 120:67:@1302.4]
  wire  _T_2758; // @[StoreQueue.scala 120:64:@1303.4]
  wire  validEntriesInLoadQ_10; // @[StoreQueue.scala 119:90:@1304.4]
  wire  _T_2762; // @[StoreQueue.scala 120:17:@1306.4]
  wire  _T_2764; // @[StoreQueue.scala 120:35:@1307.4]
  wire  _T_2765; // @[StoreQueue.scala 120:26:@1308.4]
  wire  _T_2769; // @[StoreQueue.scala 120:81:@1310.4]
  wire  _T_2771; // @[StoreQueue.scala 120:99:@1311.4]
  wire  _T_2772; // @[StoreQueue.scala 120:90:@1312.4]
  wire  _T_2774; // @[StoreQueue.scala 120:67:@1313.4]
  wire  _T_2775; // @[StoreQueue.scala 120:64:@1314.4]
  wire  validEntriesInLoadQ_11; // @[StoreQueue.scala 119:90:@1315.4]
  wire  _T_2779; // @[StoreQueue.scala 120:17:@1317.4]
  wire  _T_2781; // @[StoreQueue.scala 120:35:@1318.4]
  wire  _T_2782; // @[StoreQueue.scala 120:26:@1319.4]
  wire  _T_2786; // @[StoreQueue.scala 120:81:@1321.4]
  wire  _T_2788; // @[StoreQueue.scala 120:99:@1322.4]
  wire  _T_2789; // @[StoreQueue.scala 120:90:@1323.4]
  wire  _T_2791; // @[StoreQueue.scala 120:67:@1324.4]
  wire  _T_2792; // @[StoreQueue.scala 120:64:@1325.4]
  wire  validEntriesInLoadQ_12; // @[StoreQueue.scala 119:90:@1326.4]
  wire  _T_2796; // @[StoreQueue.scala 120:17:@1328.4]
  wire  _T_2798; // @[StoreQueue.scala 120:35:@1329.4]
  wire  _T_2799; // @[StoreQueue.scala 120:26:@1330.4]
  wire  _T_2803; // @[StoreQueue.scala 120:81:@1332.4]
  wire  _T_2805; // @[StoreQueue.scala 120:99:@1333.4]
  wire  _T_2806; // @[StoreQueue.scala 120:90:@1334.4]
  wire  _T_2808; // @[StoreQueue.scala 120:67:@1335.4]
  wire  _T_2809; // @[StoreQueue.scala 120:64:@1336.4]
  wire  validEntriesInLoadQ_13; // @[StoreQueue.scala 119:90:@1337.4]
  wire  _T_2813; // @[StoreQueue.scala 120:17:@1339.4]
  wire  _T_2815; // @[StoreQueue.scala 120:35:@1340.4]
  wire  _T_2816; // @[StoreQueue.scala 120:26:@1341.4]
  wire  _T_2820; // @[StoreQueue.scala 120:81:@1343.4]
  wire  _T_2822; // @[StoreQueue.scala 120:99:@1344.4]
  wire  _T_2823; // @[StoreQueue.scala 120:90:@1345.4]
  wire  _T_2825; // @[StoreQueue.scala 120:67:@1346.4]
  wire  _T_2826; // @[StoreQueue.scala 120:64:@1347.4]
  wire  validEntriesInLoadQ_14; // @[StoreQueue.scala 119:90:@1348.4]
  wire  validEntriesInLoadQ_15; // @[StoreQueue.scala 119:90:@1359.4]
  wire [3:0] _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  wire  _T_2869; // @[StoreQueue.scala 126:96:@1377.4]
  wire  loadsToCheck_0; // @[StoreQueue.scala 126:83:@1385.4]
  wire  _T_2899; // @[StoreQueue.scala 127:37:@1388.4]
  wire  _T_2900; // @[StoreQueue.scala 127:28:@1389.4]
  wire  _T_2905; // @[StoreQueue.scala 127:71:@1390.4]
  wire  _T_2908; // @[StoreQueue.scala 127:79:@1392.4]
  wire  _T_2910; // @[StoreQueue.scala 127:55:@1393.4]
  wire  loadsToCheck_1; // @[StoreQueue.scala 126:83:@1394.4]
  wire  _T_2922; // @[StoreQueue.scala 127:37:@1397.4]
  wire  _T_2923; // @[StoreQueue.scala 127:28:@1398.4]
  wire  _T_2928; // @[StoreQueue.scala 127:71:@1399.4]
  wire  _T_2931; // @[StoreQueue.scala 127:79:@1401.4]
  wire  _T_2933; // @[StoreQueue.scala 127:55:@1402.4]
  wire  loadsToCheck_2; // @[StoreQueue.scala 126:83:@1403.4]
  wire  _T_2945; // @[StoreQueue.scala 127:37:@1406.4]
  wire  _T_2946; // @[StoreQueue.scala 127:28:@1407.4]
  wire  _T_2951; // @[StoreQueue.scala 127:71:@1408.4]
  wire  _T_2954; // @[StoreQueue.scala 127:79:@1410.4]
  wire  _T_2956; // @[StoreQueue.scala 127:55:@1411.4]
  wire  loadsToCheck_3; // @[StoreQueue.scala 126:83:@1412.4]
  wire  _T_2968; // @[StoreQueue.scala 127:37:@1415.4]
  wire  _T_2969; // @[StoreQueue.scala 127:28:@1416.4]
  wire  _T_2974; // @[StoreQueue.scala 127:71:@1417.4]
  wire  _T_2977; // @[StoreQueue.scala 127:79:@1419.4]
  wire  _T_2979; // @[StoreQueue.scala 127:55:@1420.4]
  wire  loadsToCheck_4; // @[StoreQueue.scala 126:83:@1421.4]
  wire  _T_2991; // @[StoreQueue.scala 127:37:@1424.4]
  wire  _T_2992; // @[StoreQueue.scala 127:28:@1425.4]
  wire  _T_2997; // @[StoreQueue.scala 127:71:@1426.4]
  wire  _T_3000; // @[StoreQueue.scala 127:79:@1428.4]
  wire  _T_3002; // @[StoreQueue.scala 127:55:@1429.4]
  wire  loadsToCheck_5; // @[StoreQueue.scala 126:83:@1430.4]
  wire  _T_3014; // @[StoreQueue.scala 127:37:@1433.4]
  wire  _T_3015; // @[StoreQueue.scala 127:28:@1434.4]
  wire  _T_3020; // @[StoreQueue.scala 127:71:@1435.4]
  wire  _T_3023; // @[StoreQueue.scala 127:79:@1437.4]
  wire  _T_3025; // @[StoreQueue.scala 127:55:@1438.4]
  wire  loadsToCheck_6; // @[StoreQueue.scala 126:83:@1439.4]
  wire  _T_3037; // @[StoreQueue.scala 127:37:@1442.4]
  wire  _T_3038; // @[StoreQueue.scala 127:28:@1443.4]
  wire  _T_3043; // @[StoreQueue.scala 127:71:@1444.4]
  wire  _T_3046; // @[StoreQueue.scala 127:79:@1446.4]
  wire  _T_3048; // @[StoreQueue.scala 127:55:@1447.4]
  wire  loadsToCheck_7; // @[StoreQueue.scala 126:83:@1448.4]
  wire  _T_3060; // @[StoreQueue.scala 127:37:@1451.4]
  wire  _T_3061; // @[StoreQueue.scala 127:28:@1452.4]
  wire  _T_3066; // @[StoreQueue.scala 127:71:@1453.4]
  wire  _T_3069; // @[StoreQueue.scala 127:79:@1455.4]
  wire  _T_3071; // @[StoreQueue.scala 127:55:@1456.4]
  wire  loadsToCheck_8; // @[StoreQueue.scala 126:83:@1457.4]
  wire  _T_3083; // @[StoreQueue.scala 127:37:@1460.4]
  wire  _T_3084; // @[StoreQueue.scala 127:28:@1461.4]
  wire  _T_3089; // @[StoreQueue.scala 127:71:@1462.4]
  wire  _T_3092; // @[StoreQueue.scala 127:79:@1464.4]
  wire  _T_3094; // @[StoreQueue.scala 127:55:@1465.4]
  wire  loadsToCheck_9; // @[StoreQueue.scala 126:83:@1466.4]
  wire  _T_3106; // @[StoreQueue.scala 127:37:@1469.4]
  wire  _T_3107; // @[StoreQueue.scala 127:28:@1470.4]
  wire  _T_3112; // @[StoreQueue.scala 127:71:@1471.4]
  wire  _T_3115; // @[StoreQueue.scala 127:79:@1473.4]
  wire  _T_3117; // @[StoreQueue.scala 127:55:@1474.4]
  wire  loadsToCheck_10; // @[StoreQueue.scala 126:83:@1475.4]
  wire  _T_3129; // @[StoreQueue.scala 127:37:@1478.4]
  wire  _T_3130; // @[StoreQueue.scala 127:28:@1479.4]
  wire  _T_3135; // @[StoreQueue.scala 127:71:@1480.4]
  wire  _T_3138; // @[StoreQueue.scala 127:79:@1482.4]
  wire  _T_3140; // @[StoreQueue.scala 127:55:@1483.4]
  wire  loadsToCheck_11; // @[StoreQueue.scala 126:83:@1484.4]
  wire  _T_3152; // @[StoreQueue.scala 127:37:@1487.4]
  wire  _T_3153; // @[StoreQueue.scala 127:28:@1488.4]
  wire  _T_3158; // @[StoreQueue.scala 127:71:@1489.4]
  wire  _T_3161; // @[StoreQueue.scala 127:79:@1491.4]
  wire  _T_3163; // @[StoreQueue.scala 127:55:@1492.4]
  wire  loadsToCheck_12; // @[StoreQueue.scala 126:83:@1493.4]
  wire  _T_3175; // @[StoreQueue.scala 127:37:@1496.4]
  wire  _T_3176; // @[StoreQueue.scala 127:28:@1497.4]
  wire  _T_3181; // @[StoreQueue.scala 127:71:@1498.4]
  wire  _T_3184; // @[StoreQueue.scala 127:79:@1500.4]
  wire  _T_3186; // @[StoreQueue.scala 127:55:@1501.4]
  wire  loadsToCheck_13; // @[StoreQueue.scala 126:83:@1502.4]
  wire  _T_3198; // @[StoreQueue.scala 127:37:@1505.4]
  wire  _T_3199; // @[StoreQueue.scala 127:28:@1506.4]
  wire  _T_3204; // @[StoreQueue.scala 127:71:@1507.4]
  wire  _T_3207; // @[StoreQueue.scala 127:79:@1509.4]
  wire  _T_3209; // @[StoreQueue.scala 127:55:@1510.4]
  wire  loadsToCheck_14; // @[StoreQueue.scala 126:83:@1511.4]
  wire  _T_3221; // @[StoreQueue.scala 127:37:@1514.4]
  wire  loadsToCheck_15; // @[StoreQueue.scala 126:83:@1520.4]
  wire  _T_3255; // @[StoreQueue.scala 133:16:@1538.4]
  wire  _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  wire  entriesToCheck_0; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _T_3260; // @[StoreQueue.scala 133:16:@1540.4]
  wire  entriesToCheck_1; // @[StoreQueue.scala 133:24:@1541.4]
  wire  _T_3265; // @[StoreQueue.scala 133:16:@1542.4]
  wire  entriesToCheck_2; // @[StoreQueue.scala 133:24:@1543.4]
  wire  _T_3270; // @[StoreQueue.scala 133:16:@1544.4]
  wire  entriesToCheck_3; // @[StoreQueue.scala 133:24:@1545.4]
  wire  _T_3275; // @[StoreQueue.scala 133:16:@1546.4]
  wire  entriesToCheck_4; // @[StoreQueue.scala 133:24:@1547.4]
  wire  _T_3280; // @[StoreQueue.scala 133:16:@1548.4]
  wire  entriesToCheck_5; // @[StoreQueue.scala 133:24:@1549.4]
  wire  _T_3285; // @[StoreQueue.scala 133:16:@1550.4]
  wire  entriesToCheck_6; // @[StoreQueue.scala 133:24:@1551.4]
  wire  _T_3290; // @[StoreQueue.scala 133:16:@1552.4]
  wire  entriesToCheck_7; // @[StoreQueue.scala 133:24:@1553.4]
  wire  _T_3295; // @[StoreQueue.scala 133:16:@1554.4]
  wire  entriesToCheck_8; // @[StoreQueue.scala 133:24:@1555.4]
  wire  _T_3300; // @[StoreQueue.scala 133:16:@1556.4]
  wire  entriesToCheck_9; // @[StoreQueue.scala 133:24:@1557.4]
  wire  _T_3305; // @[StoreQueue.scala 133:16:@1558.4]
  wire  entriesToCheck_10; // @[StoreQueue.scala 133:24:@1559.4]
  wire  _T_3310; // @[StoreQueue.scala 133:16:@1560.4]
  wire  entriesToCheck_11; // @[StoreQueue.scala 133:24:@1561.4]
  wire  _T_3315; // @[StoreQueue.scala 133:16:@1562.4]
  wire  entriesToCheck_12; // @[StoreQueue.scala 133:24:@1563.4]
  wire  _T_3320; // @[StoreQueue.scala 133:16:@1564.4]
  wire  entriesToCheck_13; // @[StoreQueue.scala 133:24:@1565.4]
  wire  _T_3325; // @[StoreQueue.scala 133:16:@1566.4]
  wire  entriesToCheck_14; // @[StoreQueue.scala 133:24:@1567.4]
  wire  _T_3330; // @[StoreQueue.scala 133:16:@1568.4]
  wire  entriesToCheck_15; // @[StoreQueue.scala 133:24:@1569.4]
  wire  _T_3378; // @[StoreQueue.scala 140:34:@1588.4]
  wire  _T_3379; // @[StoreQueue.scala 140:64:@1589.4]
  wire [31:0] _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_911; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3383; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3384; // @[StoreQueue.scala 141:36:@1591.4]
  wire  noConflicts_0; // @[StoreQueue.scala 140:95:@1592.4]
  wire  _T_3387; // @[StoreQueue.scala 140:34:@1594.4]
  wire  _T_3388; // @[StoreQueue.scala 140:64:@1595.4]
  wire  _T_3392; // @[StoreQueue.scala 141:51:@1596.4]
  wire  _T_3393; // @[StoreQueue.scala 141:36:@1597.4]
  wire  noConflicts_1; // @[StoreQueue.scala 140:95:@1598.4]
  wire  _T_3396; // @[StoreQueue.scala 140:34:@1600.4]
  wire  _T_3397; // @[StoreQueue.scala 140:64:@1601.4]
  wire  _T_3401; // @[StoreQueue.scala 141:51:@1602.4]
  wire  _T_3402; // @[StoreQueue.scala 141:36:@1603.4]
  wire  noConflicts_2; // @[StoreQueue.scala 140:95:@1604.4]
  wire  _T_3405; // @[StoreQueue.scala 140:34:@1606.4]
  wire  _T_3406; // @[StoreQueue.scala 140:64:@1607.4]
  wire  _T_3410; // @[StoreQueue.scala 141:51:@1608.4]
  wire  _T_3411; // @[StoreQueue.scala 141:36:@1609.4]
  wire  noConflicts_3; // @[StoreQueue.scala 140:95:@1610.4]
  wire  _T_3414; // @[StoreQueue.scala 140:34:@1612.4]
  wire  _T_3415; // @[StoreQueue.scala 140:64:@1613.4]
  wire  _T_3419; // @[StoreQueue.scala 141:51:@1614.4]
  wire  _T_3420; // @[StoreQueue.scala 141:36:@1615.4]
  wire  noConflicts_4; // @[StoreQueue.scala 140:95:@1616.4]
  wire  _T_3423; // @[StoreQueue.scala 140:34:@1618.4]
  wire  _T_3424; // @[StoreQueue.scala 140:64:@1619.4]
  wire  _T_3428; // @[StoreQueue.scala 141:51:@1620.4]
  wire  _T_3429; // @[StoreQueue.scala 141:36:@1621.4]
  wire  noConflicts_5; // @[StoreQueue.scala 140:95:@1622.4]
  wire  _T_3432; // @[StoreQueue.scala 140:34:@1624.4]
  wire  _T_3433; // @[StoreQueue.scala 140:64:@1625.4]
  wire  _T_3437; // @[StoreQueue.scala 141:51:@1626.4]
  wire  _T_3438; // @[StoreQueue.scala 141:36:@1627.4]
  wire  noConflicts_6; // @[StoreQueue.scala 140:95:@1628.4]
  wire  _T_3441; // @[StoreQueue.scala 140:34:@1630.4]
  wire  _T_3442; // @[StoreQueue.scala 140:64:@1631.4]
  wire  _T_3446; // @[StoreQueue.scala 141:51:@1632.4]
  wire  _T_3447; // @[StoreQueue.scala 141:36:@1633.4]
  wire  noConflicts_7; // @[StoreQueue.scala 140:95:@1634.4]
  wire  _T_3450; // @[StoreQueue.scala 140:34:@1636.4]
  wire  _T_3451; // @[StoreQueue.scala 140:64:@1637.4]
  wire  _T_3455; // @[StoreQueue.scala 141:51:@1638.4]
  wire  _T_3456; // @[StoreQueue.scala 141:36:@1639.4]
  wire  noConflicts_8; // @[StoreQueue.scala 140:95:@1640.4]
  wire  _T_3459; // @[StoreQueue.scala 140:34:@1642.4]
  wire  _T_3460; // @[StoreQueue.scala 140:64:@1643.4]
  wire  _T_3464; // @[StoreQueue.scala 141:51:@1644.4]
  wire  _T_3465; // @[StoreQueue.scala 141:36:@1645.4]
  wire  noConflicts_9; // @[StoreQueue.scala 140:95:@1646.4]
  wire  _T_3468; // @[StoreQueue.scala 140:34:@1648.4]
  wire  _T_3469; // @[StoreQueue.scala 140:64:@1649.4]
  wire  _T_3473; // @[StoreQueue.scala 141:51:@1650.4]
  wire  _T_3474; // @[StoreQueue.scala 141:36:@1651.4]
  wire  noConflicts_10; // @[StoreQueue.scala 140:95:@1652.4]
  wire  _T_3477; // @[StoreQueue.scala 140:34:@1654.4]
  wire  _T_3478; // @[StoreQueue.scala 140:64:@1655.4]
  wire  _T_3482; // @[StoreQueue.scala 141:51:@1656.4]
  wire  _T_3483; // @[StoreQueue.scala 141:36:@1657.4]
  wire  noConflicts_11; // @[StoreQueue.scala 140:95:@1658.4]
  wire  _T_3486; // @[StoreQueue.scala 140:34:@1660.4]
  wire  _T_3487; // @[StoreQueue.scala 140:64:@1661.4]
  wire  _T_3491; // @[StoreQueue.scala 141:51:@1662.4]
  wire  _T_3492; // @[StoreQueue.scala 141:36:@1663.4]
  wire  noConflicts_12; // @[StoreQueue.scala 140:95:@1664.4]
  wire  _T_3495; // @[StoreQueue.scala 140:34:@1666.4]
  wire  _T_3496; // @[StoreQueue.scala 140:64:@1667.4]
  wire  _T_3500; // @[StoreQueue.scala 141:51:@1668.4]
  wire  _T_3501; // @[StoreQueue.scala 141:36:@1669.4]
  wire  noConflicts_13; // @[StoreQueue.scala 140:95:@1670.4]
  wire  _T_3504; // @[StoreQueue.scala 140:34:@1672.4]
  wire  _T_3505; // @[StoreQueue.scala 140:64:@1673.4]
  wire  _T_3509; // @[StoreQueue.scala 141:51:@1674.4]
  wire  _T_3510; // @[StoreQueue.scala 141:36:@1675.4]
  wire  noConflicts_14; // @[StoreQueue.scala 140:95:@1676.4]
  wire  _T_3513; // @[StoreQueue.scala 140:34:@1678.4]
  wire  _T_3514; // @[StoreQueue.scala 140:64:@1679.4]
  wire  _T_3518; // @[StoreQueue.scala 141:51:@1680.4]
  wire  _T_3519; // @[StoreQueue.scala 141:36:@1681.4]
  wire  noConflicts_15; // @[StoreQueue.scala 140:95:@1682.4]
  wire  _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_927; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _T_3527; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_959; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3532; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3533; // @[StoreQueue.scala 154:63:@1686.4]
  wire  _T_3536; // @[StoreQueue.scala 154:109:@1688.4]
  wire  _T_3537; // @[StoreQueue.scala 154:109:@1689.4]
  wire  _T_3538; // @[StoreQueue.scala 154:109:@1690.4]
  wire  _T_3539; // @[StoreQueue.scala 154:109:@1691.4]
  wire  _T_3540; // @[StoreQueue.scala 154:109:@1692.4]
  wire  _T_3541; // @[StoreQueue.scala 154:109:@1693.4]
  wire  _T_3542; // @[StoreQueue.scala 154:109:@1694.4]
  wire  _T_3543; // @[StoreQueue.scala 154:109:@1695.4]
  wire  _T_3544; // @[StoreQueue.scala 154:109:@1696.4]
  wire  _T_3545; // @[StoreQueue.scala 154:109:@1697.4]
  wire  _T_3546; // @[StoreQueue.scala 154:109:@1698.4]
  wire  _T_3547; // @[StoreQueue.scala 154:109:@1699.4]
  wire  _T_3548; // @[StoreQueue.scala 154:109:@1700.4]
  wire  _T_3549; // @[StoreQueue.scala 154:109:@1701.4]
  wire  _T_3550; // @[StoreQueue.scala 154:109:@1702.4]
  wire  storeRequest; // @[StoreQueue.scala 154:88:@1703.4]
  wire  _T_3553; // @[StoreQueue.scala 164:23:@1708.6]
  wire  _T_3554; // @[StoreQueue.scala 164:43:@1709.6]
  wire  _T_3555; // @[StoreQueue.scala 164:59:@1710.6]
  wire  _GEN_960; // @[StoreQueue.scala 164:86:@1711.6]
  wire  _GEN_961; // @[StoreQueue.scala 162:37:@1704.4]
  wire  _T_3559; // @[StoreQueue.scala 164:23:@1718.6]
  wire  _T_3560; // @[StoreQueue.scala 164:43:@1719.6]
  wire  _T_3561; // @[StoreQueue.scala 164:59:@1720.6]
  wire  _GEN_962; // @[StoreQueue.scala 164:86:@1721.6]
  wire  _GEN_963; // @[StoreQueue.scala 162:37:@1714.4]
  wire  _T_3565; // @[StoreQueue.scala 164:23:@1728.6]
  wire  _T_3566; // @[StoreQueue.scala 164:43:@1729.6]
  wire  _T_3567; // @[StoreQueue.scala 164:59:@1730.6]
  wire  _GEN_964; // @[StoreQueue.scala 164:86:@1731.6]
  wire  _GEN_965; // @[StoreQueue.scala 162:37:@1724.4]
  wire  _T_3571; // @[StoreQueue.scala 164:23:@1738.6]
  wire  _T_3572; // @[StoreQueue.scala 164:43:@1739.6]
  wire  _T_3573; // @[StoreQueue.scala 164:59:@1740.6]
  wire  _GEN_966; // @[StoreQueue.scala 164:86:@1741.6]
  wire  _GEN_967; // @[StoreQueue.scala 162:37:@1734.4]
  wire  _T_3577; // @[StoreQueue.scala 164:23:@1748.6]
  wire  _T_3578; // @[StoreQueue.scala 164:43:@1749.6]
  wire  _T_3579; // @[StoreQueue.scala 164:59:@1750.6]
  wire  _GEN_968; // @[StoreQueue.scala 164:86:@1751.6]
  wire  _GEN_969; // @[StoreQueue.scala 162:37:@1744.4]
  wire  _T_3583; // @[StoreQueue.scala 164:23:@1758.6]
  wire  _T_3584; // @[StoreQueue.scala 164:43:@1759.6]
  wire  _T_3585; // @[StoreQueue.scala 164:59:@1760.6]
  wire  _GEN_970; // @[StoreQueue.scala 164:86:@1761.6]
  wire  _GEN_971; // @[StoreQueue.scala 162:37:@1754.4]
  wire  _T_3589; // @[StoreQueue.scala 164:23:@1768.6]
  wire  _T_3590; // @[StoreQueue.scala 164:43:@1769.6]
  wire  _T_3591; // @[StoreQueue.scala 164:59:@1770.6]
  wire  _GEN_972; // @[StoreQueue.scala 164:86:@1771.6]
  wire  _GEN_973; // @[StoreQueue.scala 162:37:@1764.4]
  wire  _T_3595; // @[StoreQueue.scala 164:23:@1778.6]
  wire  _T_3596; // @[StoreQueue.scala 164:43:@1779.6]
  wire  _T_3597; // @[StoreQueue.scala 164:59:@1780.6]
  wire  _GEN_974; // @[StoreQueue.scala 164:86:@1781.6]
  wire  _GEN_975; // @[StoreQueue.scala 162:37:@1774.4]
  wire  _T_3601; // @[StoreQueue.scala 164:23:@1788.6]
  wire  _T_3602; // @[StoreQueue.scala 164:43:@1789.6]
  wire  _T_3603; // @[StoreQueue.scala 164:59:@1790.6]
  wire  _GEN_976; // @[StoreQueue.scala 164:86:@1791.6]
  wire  _GEN_977; // @[StoreQueue.scala 162:37:@1784.4]
  wire  _T_3607; // @[StoreQueue.scala 164:23:@1798.6]
  wire  _T_3608; // @[StoreQueue.scala 164:43:@1799.6]
  wire  _T_3609; // @[StoreQueue.scala 164:59:@1800.6]
  wire  _GEN_978; // @[StoreQueue.scala 164:86:@1801.6]
  wire  _GEN_979; // @[StoreQueue.scala 162:37:@1794.4]
  wire  _T_3613; // @[StoreQueue.scala 164:23:@1808.6]
  wire  _T_3614; // @[StoreQueue.scala 164:43:@1809.6]
  wire  _T_3615; // @[StoreQueue.scala 164:59:@1810.6]
  wire  _GEN_980; // @[StoreQueue.scala 164:86:@1811.6]
  wire  _GEN_981; // @[StoreQueue.scala 162:37:@1804.4]
  wire  _T_3619; // @[StoreQueue.scala 164:23:@1818.6]
  wire  _T_3620; // @[StoreQueue.scala 164:43:@1819.6]
  wire  _T_3621; // @[StoreQueue.scala 164:59:@1820.6]
  wire  _GEN_982; // @[StoreQueue.scala 164:86:@1821.6]
  wire  _GEN_983; // @[StoreQueue.scala 162:37:@1814.4]
  wire  _T_3625; // @[StoreQueue.scala 164:23:@1828.6]
  wire  _T_3626; // @[StoreQueue.scala 164:43:@1829.6]
  wire  _T_3627; // @[StoreQueue.scala 164:59:@1830.6]
  wire  _GEN_984; // @[StoreQueue.scala 164:86:@1831.6]
  wire  _GEN_985; // @[StoreQueue.scala 162:37:@1824.4]
  wire  _T_3631; // @[StoreQueue.scala 164:23:@1838.6]
  wire  _T_3632; // @[StoreQueue.scala 164:43:@1839.6]
  wire  _T_3633; // @[StoreQueue.scala 164:59:@1840.6]
  wire  _GEN_986; // @[StoreQueue.scala 164:86:@1841.6]
  wire  _GEN_987; // @[StoreQueue.scala 162:37:@1834.4]
  wire  _T_3637; // @[StoreQueue.scala 164:23:@1848.6]
  wire  _T_3638; // @[StoreQueue.scala 164:43:@1849.6]
  wire  _T_3639; // @[StoreQueue.scala 164:59:@1850.6]
  wire  _GEN_988; // @[StoreQueue.scala 164:86:@1851.6]
  wire  _GEN_989; // @[StoreQueue.scala 162:37:@1844.4]
  wire  _T_3643; // @[StoreQueue.scala 164:23:@1858.6]
  wire  _T_3644; // @[StoreQueue.scala 164:43:@1859.6]
  wire  _T_3645; // @[StoreQueue.scala 164:59:@1860.6]
  wire  _GEN_990; // @[StoreQueue.scala 164:86:@1861.6]
  wire  _GEN_991; // @[StoreQueue.scala 162:37:@1854.4]
  wire  entriesPorts_0_0; // @[StoreQueue.scala 180:72:@1865.4]
  wire  entriesPorts_0_1; // @[StoreQueue.scala 180:72:@1867.4]
  wire  entriesPorts_0_2; // @[StoreQueue.scala 180:72:@1869.4]
  wire  entriesPorts_0_3; // @[StoreQueue.scala 180:72:@1871.4]
  wire  entriesPorts_0_4; // @[StoreQueue.scala 180:72:@1873.4]
  wire  entriesPorts_0_5; // @[StoreQueue.scala 180:72:@1875.4]
  wire  entriesPorts_0_6; // @[StoreQueue.scala 180:72:@1877.4]
  wire  entriesPorts_0_7; // @[StoreQueue.scala 180:72:@1879.4]
  wire  entriesPorts_0_8; // @[StoreQueue.scala 180:72:@1881.4]
  wire  entriesPorts_0_9; // @[StoreQueue.scala 180:72:@1883.4]
  wire  entriesPorts_0_10; // @[StoreQueue.scala 180:72:@1885.4]
  wire  entriesPorts_0_11; // @[StoreQueue.scala 180:72:@1887.4]
  wire  entriesPorts_0_12; // @[StoreQueue.scala 180:72:@1889.4]
  wire  entriesPorts_0_13; // @[StoreQueue.scala 180:72:@1891.4]
  wire  entriesPorts_0_14; // @[StoreQueue.scala 180:72:@1893.4]
  wire  entriesPorts_0_15; // @[StoreQueue.scala 180:72:@1895.4]
  wire  _T_4378; // @[StoreQueue.scala 192:91:@1931.4]
  wire  _T_4379; // @[StoreQueue.scala 192:88:@1932.4]
  wire  _T_4381; // @[StoreQueue.scala 192:91:@1933.4]
  wire  _T_4382; // @[StoreQueue.scala 192:88:@1934.4]
  wire  _T_4384; // @[StoreQueue.scala 192:91:@1935.4]
  wire  _T_4385; // @[StoreQueue.scala 192:88:@1936.4]
  wire  _T_4387; // @[StoreQueue.scala 192:91:@1937.4]
  wire  _T_4388; // @[StoreQueue.scala 192:88:@1938.4]
  wire  _T_4390; // @[StoreQueue.scala 192:91:@1939.4]
  wire  _T_4391; // @[StoreQueue.scala 192:88:@1940.4]
  wire  _T_4393; // @[StoreQueue.scala 192:91:@1941.4]
  wire  _T_4394; // @[StoreQueue.scala 192:88:@1942.4]
  wire  _T_4396; // @[StoreQueue.scala 192:91:@1943.4]
  wire  _T_4397; // @[StoreQueue.scala 192:88:@1944.4]
  wire  _T_4399; // @[StoreQueue.scala 192:91:@1945.4]
  wire  _T_4400; // @[StoreQueue.scala 192:88:@1946.4]
  wire  _T_4402; // @[StoreQueue.scala 192:91:@1947.4]
  wire  _T_4403; // @[StoreQueue.scala 192:88:@1948.4]
  wire  _T_4405; // @[StoreQueue.scala 192:91:@1949.4]
  wire  _T_4406; // @[StoreQueue.scala 192:88:@1950.4]
  wire  _T_4408; // @[StoreQueue.scala 192:91:@1951.4]
  wire  _T_4409; // @[StoreQueue.scala 192:88:@1952.4]
  wire  _T_4411; // @[StoreQueue.scala 192:91:@1953.4]
  wire  _T_4412; // @[StoreQueue.scala 192:88:@1954.4]
  wire  _T_4414; // @[StoreQueue.scala 192:91:@1955.4]
  wire  _T_4415; // @[StoreQueue.scala 192:88:@1956.4]
  wire  _T_4417; // @[StoreQueue.scala 192:91:@1957.4]
  wire  _T_4418; // @[StoreQueue.scala 192:88:@1958.4]
  wire  _T_4420; // @[StoreQueue.scala 192:91:@1959.4]
  wire  _T_4421; // @[StoreQueue.scala 192:88:@1960.4]
  wire  _T_4423; // @[StoreQueue.scala 192:91:@1961.4]
  wire  _T_4424; // @[StoreQueue.scala 192:88:@1962.4]
  wire  _T_4448; // @[StoreQueue.scala 193:91:@1980.4]
  wire  _T_4449; // @[StoreQueue.scala 193:88:@1981.4]
  wire  _T_4451; // @[StoreQueue.scala 193:91:@1982.4]
  wire  _T_4452; // @[StoreQueue.scala 193:88:@1983.4]
  wire  _T_4454; // @[StoreQueue.scala 193:91:@1984.4]
  wire  _T_4455; // @[StoreQueue.scala 193:88:@1985.4]
  wire  _T_4457; // @[StoreQueue.scala 193:91:@1986.4]
  wire  _T_4458; // @[StoreQueue.scala 193:88:@1987.4]
  wire  _T_4460; // @[StoreQueue.scala 193:91:@1988.4]
  wire  _T_4461; // @[StoreQueue.scala 193:88:@1989.4]
  wire  _T_4463; // @[StoreQueue.scala 193:91:@1990.4]
  wire  _T_4464; // @[StoreQueue.scala 193:88:@1991.4]
  wire  _T_4466; // @[StoreQueue.scala 193:91:@1992.4]
  wire  _T_4467; // @[StoreQueue.scala 193:88:@1993.4]
  wire  _T_4469; // @[StoreQueue.scala 193:91:@1994.4]
  wire  _T_4470; // @[StoreQueue.scala 193:88:@1995.4]
  wire  _T_4472; // @[StoreQueue.scala 193:91:@1996.4]
  wire  _T_4473; // @[StoreQueue.scala 193:88:@1997.4]
  wire  _T_4475; // @[StoreQueue.scala 193:91:@1998.4]
  wire  _T_4476; // @[StoreQueue.scala 193:88:@1999.4]
  wire  _T_4478; // @[StoreQueue.scala 193:91:@2000.4]
  wire  _T_4479; // @[StoreQueue.scala 193:88:@2001.4]
  wire  _T_4481; // @[StoreQueue.scala 193:91:@2002.4]
  wire  _T_4482; // @[StoreQueue.scala 193:88:@2003.4]
  wire  _T_4484; // @[StoreQueue.scala 193:91:@2004.4]
  wire  _T_4485; // @[StoreQueue.scala 193:88:@2005.4]
  wire  _T_4487; // @[StoreQueue.scala 193:91:@2006.4]
  wire  _T_4488; // @[StoreQueue.scala 193:88:@2007.4]
  wire  _T_4490; // @[StoreQueue.scala 193:91:@2008.4]
  wire  _T_4491; // @[StoreQueue.scala 193:88:@2009.4]
  wire  _T_4493; // @[StoreQueue.scala 193:91:@2010.4]
  wire  _T_4494; // @[StoreQueue.scala 193:88:@2011.4]
  wire [15:0] _T_4519; // @[OneHot.scala 52:12:@2030.4]
  wire  _T_4521; // @[util.scala 33:60:@2032.4]
  wire  _T_4522; // @[util.scala 33:60:@2033.4]
  wire  _T_4523; // @[util.scala 33:60:@2034.4]
  wire  _T_4524; // @[util.scala 33:60:@2035.4]
  wire  _T_4525; // @[util.scala 33:60:@2036.4]
  wire  _T_4526; // @[util.scala 33:60:@2037.4]
  wire  _T_4527; // @[util.scala 33:60:@2038.4]
  wire  _T_4528; // @[util.scala 33:60:@2039.4]
  wire  _T_4529; // @[util.scala 33:60:@2040.4]
  wire  _T_4530; // @[util.scala 33:60:@2041.4]
  wire  _T_4531; // @[util.scala 33:60:@2042.4]
  wire  _T_4532; // @[util.scala 33:60:@2043.4]
  wire  _T_4533; // @[util.scala 33:60:@2044.4]
  wire  _T_4534; // @[util.scala 33:60:@2045.4]
  wire  _T_4535; // @[util.scala 33:60:@2046.4]
  wire  _T_4536; // @[util.scala 33:60:@2047.4]
  wire [15:0] _T_4577; // @[Mux.scala 31:69:@2065.4]
  wire [15:0] _T_4578; // @[Mux.scala 31:69:@2066.4]
  wire [15:0] _T_4579; // @[Mux.scala 31:69:@2067.4]
  wire [15:0] _T_4580; // @[Mux.scala 31:69:@2068.4]
  wire [15:0] _T_4581; // @[Mux.scala 31:69:@2069.4]
  wire [15:0] _T_4582; // @[Mux.scala 31:69:@2070.4]
  wire [15:0] _T_4583; // @[Mux.scala 31:69:@2071.4]
  wire [15:0] _T_4584; // @[Mux.scala 31:69:@2072.4]
  wire [15:0] _T_4585; // @[Mux.scala 31:69:@2073.4]
  wire [15:0] _T_4586; // @[Mux.scala 31:69:@2074.4]
  wire [15:0] _T_4587; // @[Mux.scala 31:69:@2075.4]
  wire [15:0] _T_4588; // @[Mux.scala 31:69:@2076.4]
  wire [15:0] _T_4589; // @[Mux.scala 31:69:@2077.4]
  wire [15:0] _T_4590; // @[Mux.scala 31:69:@2078.4]
  wire [15:0] _T_4591; // @[Mux.scala 31:69:@2079.4]
  wire [15:0] _T_4592; // @[Mux.scala 31:69:@2080.4]
  wire  _T_4593; // @[OneHot.scala 66:30:@2081.4]
  wire  _T_4594; // @[OneHot.scala 66:30:@2082.4]
  wire  _T_4595; // @[OneHot.scala 66:30:@2083.4]
  wire  _T_4596; // @[OneHot.scala 66:30:@2084.4]
  wire  _T_4597; // @[OneHot.scala 66:30:@2085.4]
  wire  _T_4598; // @[OneHot.scala 66:30:@2086.4]
  wire  _T_4599; // @[OneHot.scala 66:30:@2087.4]
  wire  _T_4600; // @[OneHot.scala 66:30:@2088.4]
  wire  _T_4601; // @[OneHot.scala 66:30:@2089.4]
  wire  _T_4602; // @[OneHot.scala 66:30:@2090.4]
  wire  _T_4603; // @[OneHot.scala 66:30:@2091.4]
  wire  _T_4604; // @[OneHot.scala 66:30:@2092.4]
  wire  _T_4605; // @[OneHot.scala 66:30:@2093.4]
  wire  _T_4606; // @[OneHot.scala 66:30:@2094.4]
  wire  _T_4607; // @[OneHot.scala 66:30:@2095.4]
  wire  _T_4608; // @[OneHot.scala 66:30:@2096.4]
  wire [15:0] _T_4649; // @[Mux.scala 31:69:@2114.4]
  wire [15:0] _T_4650; // @[Mux.scala 31:69:@2115.4]
  wire [15:0] _T_4651; // @[Mux.scala 31:69:@2116.4]
  wire [15:0] _T_4652; // @[Mux.scala 31:69:@2117.4]
  wire [15:0] _T_4653; // @[Mux.scala 31:69:@2118.4]
  wire [15:0] _T_4654; // @[Mux.scala 31:69:@2119.4]
  wire [15:0] _T_4655; // @[Mux.scala 31:69:@2120.4]
  wire [15:0] _T_4656; // @[Mux.scala 31:69:@2121.4]
  wire [15:0] _T_4657; // @[Mux.scala 31:69:@2122.4]
  wire [15:0] _T_4658; // @[Mux.scala 31:69:@2123.4]
  wire [15:0] _T_4659; // @[Mux.scala 31:69:@2124.4]
  wire [15:0] _T_4660; // @[Mux.scala 31:69:@2125.4]
  wire [15:0] _T_4661; // @[Mux.scala 31:69:@2126.4]
  wire [15:0] _T_4662; // @[Mux.scala 31:69:@2127.4]
  wire [15:0] _T_4663; // @[Mux.scala 31:69:@2128.4]
  wire [15:0] _T_4664; // @[Mux.scala 31:69:@2129.4]
  wire  _T_4665; // @[OneHot.scala 66:30:@2130.4]
  wire  _T_4666; // @[OneHot.scala 66:30:@2131.4]
  wire  _T_4667; // @[OneHot.scala 66:30:@2132.4]
  wire  _T_4668; // @[OneHot.scala 66:30:@2133.4]
  wire  _T_4669; // @[OneHot.scala 66:30:@2134.4]
  wire  _T_4670; // @[OneHot.scala 66:30:@2135.4]
  wire  _T_4671; // @[OneHot.scala 66:30:@2136.4]
  wire  _T_4672; // @[OneHot.scala 66:30:@2137.4]
  wire  _T_4673; // @[OneHot.scala 66:30:@2138.4]
  wire  _T_4674; // @[OneHot.scala 66:30:@2139.4]
  wire  _T_4675; // @[OneHot.scala 66:30:@2140.4]
  wire  _T_4676; // @[OneHot.scala 66:30:@2141.4]
  wire  _T_4677; // @[OneHot.scala 66:30:@2142.4]
  wire  _T_4678; // @[OneHot.scala 66:30:@2143.4]
  wire  _T_4679; // @[OneHot.scala 66:30:@2144.4]
  wire  _T_4680; // @[OneHot.scala 66:30:@2145.4]
  wire [15:0] _T_4721; // @[Mux.scala 31:69:@2163.4]
  wire [15:0] _T_4722; // @[Mux.scala 31:69:@2164.4]
  wire [15:0] _T_4723; // @[Mux.scala 31:69:@2165.4]
  wire [15:0] _T_4724; // @[Mux.scala 31:69:@2166.4]
  wire [15:0] _T_4725; // @[Mux.scala 31:69:@2167.4]
  wire [15:0] _T_4726; // @[Mux.scala 31:69:@2168.4]
  wire [15:0] _T_4727; // @[Mux.scala 31:69:@2169.4]
  wire [15:0] _T_4728; // @[Mux.scala 31:69:@2170.4]
  wire [15:0] _T_4729; // @[Mux.scala 31:69:@2171.4]
  wire [15:0] _T_4730; // @[Mux.scala 31:69:@2172.4]
  wire [15:0] _T_4731; // @[Mux.scala 31:69:@2173.4]
  wire [15:0] _T_4732; // @[Mux.scala 31:69:@2174.4]
  wire [15:0] _T_4733; // @[Mux.scala 31:69:@2175.4]
  wire [15:0] _T_4734; // @[Mux.scala 31:69:@2176.4]
  wire [15:0] _T_4735; // @[Mux.scala 31:69:@2177.4]
  wire [15:0] _T_4736; // @[Mux.scala 31:69:@2178.4]
  wire  _T_4737; // @[OneHot.scala 66:30:@2179.4]
  wire  _T_4738; // @[OneHot.scala 66:30:@2180.4]
  wire  _T_4739; // @[OneHot.scala 66:30:@2181.4]
  wire  _T_4740; // @[OneHot.scala 66:30:@2182.4]
  wire  _T_4741; // @[OneHot.scala 66:30:@2183.4]
  wire  _T_4742; // @[OneHot.scala 66:30:@2184.4]
  wire  _T_4743; // @[OneHot.scala 66:30:@2185.4]
  wire  _T_4744; // @[OneHot.scala 66:30:@2186.4]
  wire  _T_4745; // @[OneHot.scala 66:30:@2187.4]
  wire  _T_4746; // @[OneHot.scala 66:30:@2188.4]
  wire  _T_4747; // @[OneHot.scala 66:30:@2189.4]
  wire  _T_4748; // @[OneHot.scala 66:30:@2190.4]
  wire  _T_4749; // @[OneHot.scala 66:30:@2191.4]
  wire  _T_4750; // @[OneHot.scala 66:30:@2192.4]
  wire  _T_4751; // @[OneHot.scala 66:30:@2193.4]
  wire  _T_4752; // @[OneHot.scala 66:30:@2194.4]
  wire [15:0] _T_4793; // @[Mux.scala 31:69:@2212.4]
  wire [15:0] _T_4794; // @[Mux.scala 31:69:@2213.4]
  wire [15:0] _T_4795; // @[Mux.scala 31:69:@2214.4]
  wire [15:0] _T_4796; // @[Mux.scala 31:69:@2215.4]
  wire [15:0] _T_4797; // @[Mux.scala 31:69:@2216.4]
  wire [15:0] _T_4798; // @[Mux.scala 31:69:@2217.4]
  wire [15:0] _T_4799; // @[Mux.scala 31:69:@2218.4]
  wire [15:0] _T_4800; // @[Mux.scala 31:69:@2219.4]
  wire [15:0] _T_4801; // @[Mux.scala 31:69:@2220.4]
  wire [15:0] _T_4802; // @[Mux.scala 31:69:@2221.4]
  wire [15:0] _T_4803; // @[Mux.scala 31:69:@2222.4]
  wire [15:0] _T_4804; // @[Mux.scala 31:69:@2223.4]
  wire [15:0] _T_4805; // @[Mux.scala 31:69:@2224.4]
  wire [15:0] _T_4806; // @[Mux.scala 31:69:@2225.4]
  wire [15:0] _T_4807; // @[Mux.scala 31:69:@2226.4]
  wire [15:0] _T_4808; // @[Mux.scala 31:69:@2227.4]
  wire  _T_4809; // @[OneHot.scala 66:30:@2228.4]
  wire  _T_4810; // @[OneHot.scala 66:30:@2229.4]
  wire  _T_4811; // @[OneHot.scala 66:30:@2230.4]
  wire  _T_4812; // @[OneHot.scala 66:30:@2231.4]
  wire  _T_4813; // @[OneHot.scala 66:30:@2232.4]
  wire  _T_4814; // @[OneHot.scala 66:30:@2233.4]
  wire  _T_4815; // @[OneHot.scala 66:30:@2234.4]
  wire  _T_4816; // @[OneHot.scala 66:30:@2235.4]
  wire  _T_4817; // @[OneHot.scala 66:30:@2236.4]
  wire  _T_4818; // @[OneHot.scala 66:30:@2237.4]
  wire  _T_4819; // @[OneHot.scala 66:30:@2238.4]
  wire  _T_4820; // @[OneHot.scala 66:30:@2239.4]
  wire  _T_4821; // @[OneHot.scala 66:30:@2240.4]
  wire  _T_4822; // @[OneHot.scala 66:30:@2241.4]
  wire  _T_4823; // @[OneHot.scala 66:30:@2242.4]
  wire  _T_4824; // @[OneHot.scala 66:30:@2243.4]
  wire [15:0] _T_4865; // @[Mux.scala 31:69:@2261.4]
  wire [15:0] _T_4866; // @[Mux.scala 31:69:@2262.4]
  wire [15:0] _T_4867; // @[Mux.scala 31:69:@2263.4]
  wire [15:0] _T_4868; // @[Mux.scala 31:69:@2264.4]
  wire [15:0] _T_4869; // @[Mux.scala 31:69:@2265.4]
  wire [15:0] _T_4870; // @[Mux.scala 31:69:@2266.4]
  wire [15:0] _T_4871; // @[Mux.scala 31:69:@2267.4]
  wire [15:0] _T_4872; // @[Mux.scala 31:69:@2268.4]
  wire [15:0] _T_4873; // @[Mux.scala 31:69:@2269.4]
  wire [15:0] _T_4874; // @[Mux.scala 31:69:@2270.4]
  wire [15:0] _T_4875; // @[Mux.scala 31:69:@2271.4]
  wire [15:0] _T_4876; // @[Mux.scala 31:69:@2272.4]
  wire [15:0] _T_4877; // @[Mux.scala 31:69:@2273.4]
  wire [15:0] _T_4878; // @[Mux.scala 31:69:@2274.4]
  wire [15:0] _T_4879; // @[Mux.scala 31:69:@2275.4]
  wire [15:0] _T_4880; // @[Mux.scala 31:69:@2276.4]
  wire  _T_4881; // @[OneHot.scala 66:30:@2277.4]
  wire  _T_4882; // @[OneHot.scala 66:30:@2278.4]
  wire  _T_4883; // @[OneHot.scala 66:30:@2279.4]
  wire  _T_4884; // @[OneHot.scala 66:30:@2280.4]
  wire  _T_4885; // @[OneHot.scala 66:30:@2281.4]
  wire  _T_4886; // @[OneHot.scala 66:30:@2282.4]
  wire  _T_4887; // @[OneHot.scala 66:30:@2283.4]
  wire  _T_4888; // @[OneHot.scala 66:30:@2284.4]
  wire  _T_4889; // @[OneHot.scala 66:30:@2285.4]
  wire  _T_4890; // @[OneHot.scala 66:30:@2286.4]
  wire  _T_4891; // @[OneHot.scala 66:30:@2287.4]
  wire  _T_4892; // @[OneHot.scala 66:30:@2288.4]
  wire  _T_4893; // @[OneHot.scala 66:30:@2289.4]
  wire  _T_4894; // @[OneHot.scala 66:30:@2290.4]
  wire  _T_4895; // @[OneHot.scala 66:30:@2291.4]
  wire  _T_4896; // @[OneHot.scala 66:30:@2292.4]
  wire [15:0] _T_4937; // @[Mux.scala 31:69:@2310.4]
  wire [15:0] _T_4938; // @[Mux.scala 31:69:@2311.4]
  wire [15:0] _T_4939; // @[Mux.scala 31:69:@2312.4]
  wire [15:0] _T_4940; // @[Mux.scala 31:69:@2313.4]
  wire [15:0] _T_4941; // @[Mux.scala 31:69:@2314.4]
  wire [15:0] _T_4942; // @[Mux.scala 31:69:@2315.4]
  wire [15:0] _T_4943; // @[Mux.scala 31:69:@2316.4]
  wire [15:0] _T_4944; // @[Mux.scala 31:69:@2317.4]
  wire [15:0] _T_4945; // @[Mux.scala 31:69:@2318.4]
  wire [15:0] _T_4946; // @[Mux.scala 31:69:@2319.4]
  wire [15:0] _T_4947; // @[Mux.scala 31:69:@2320.4]
  wire [15:0] _T_4948; // @[Mux.scala 31:69:@2321.4]
  wire [15:0] _T_4949; // @[Mux.scala 31:69:@2322.4]
  wire [15:0] _T_4950; // @[Mux.scala 31:69:@2323.4]
  wire [15:0] _T_4951; // @[Mux.scala 31:69:@2324.4]
  wire [15:0] _T_4952; // @[Mux.scala 31:69:@2325.4]
  wire  _T_4953; // @[OneHot.scala 66:30:@2326.4]
  wire  _T_4954; // @[OneHot.scala 66:30:@2327.4]
  wire  _T_4955; // @[OneHot.scala 66:30:@2328.4]
  wire  _T_4956; // @[OneHot.scala 66:30:@2329.4]
  wire  _T_4957; // @[OneHot.scala 66:30:@2330.4]
  wire  _T_4958; // @[OneHot.scala 66:30:@2331.4]
  wire  _T_4959; // @[OneHot.scala 66:30:@2332.4]
  wire  _T_4960; // @[OneHot.scala 66:30:@2333.4]
  wire  _T_4961; // @[OneHot.scala 66:30:@2334.4]
  wire  _T_4962; // @[OneHot.scala 66:30:@2335.4]
  wire  _T_4963; // @[OneHot.scala 66:30:@2336.4]
  wire  _T_4964; // @[OneHot.scala 66:30:@2337.4]
  wire  _T_4965; // @[OneHot.scala 66:30:@2338.4]
  wire  _T_4966; // @[OneHot.scala 66:30:@2339.4]
  wire  _T_4967; // @[OneHot.scala 66:30:@2340.4]
  wire  _T_4968; // @[OneHot.scala 66:30:@2341.4]
  wire [15:0] _T_5009; // @[Mux.scala 31:69:@2359.4]
  wire [15:0] _T_5010; // @[Mux.scala 31:69:@2360.4]
  wire [15:0] _T_5011; // @[Mux.scala 31:69:@2361.4]
  wire [15:0] _T_5012; // @[Mux.scala 31:69:@2362.4]
  wire [15:0] _T_5013; // @[Mux.scala 31:69:@2363.4]
  wire [15:0] _T_5014; // @[Mux.scala 31:69:@2364.4]
  wire [15:0] _T_5015; // @[Mux.scala 31:69:@2365.4]
  wire [15:0] _T_5016; // @[Mux.scala 31:69:@2366.4]
  wire [15:0] _T_5017; // @[Mux.scala 31:69:@2367.4]
  wire [15:0] _T_5018; // @[Mux.scala 31:69:@2368.4]
  wire [15:0] _T_5019; // @[Mux.scala 31:69:@2369.4]
  wire [15:0] _T_5020; // @[Mux.scala 31:69:@2370.4]
  wire [15:0] _T_5021; // @[Mux.scala 31:69:@2371.4]
  wire [15:0] _T_5022; // @[Mux.scala 31:69:@2372.4]
  wire [15:0] _T_5023; // @[Mux.scala 31:69:@2373.4]
  wire [15:0] _T_5024; // @[Mux.scala 31:69:@2374.4]
  wire  _T_5025; // @[OneHot.scala 66:30:@2375.4]
  wire  _T_5026; // @[OneHot.scala 66:30:@2376.4]
  wire  _T_5027; // @[OneHot.scala 66:30:@2377.4]
  wire  _T_5028; // @[OneHot.scala 66:30:@2378.4]
  wire  _T_5029; // @[OneHot.scala 66:30:@2379.4]
  wire  _T_5030; // @[OneHot.scala 66:30:@2380.4]
  wire  _T_5031; // @[OneHot.scala 66:30:@2381.4]
  wire  _T_5032; // @[OneHot.scala 66:30:@2382.4]
  wire  _T_5033; // @[OneHot.scala 66:30:@2383.4]
  wire  _T_5034; // @[OneHot.scala 66:30:@2384.4]
  wire  _T_5035; // @[OneHot.scala 66:30:@2385.4]
  wire  _T_5036; // @[OneHot.scala 66:30:@2386.4]
  wire  _T_5037; // @[OneHot.scala 66:30:@2387.4]
  wire  _T_5038; // @[OneHot.scala 66:30:@2388.4]
  wire  _T_5039; // @[OneHot.scala 66:30:@2389.4]
  wire  _T_5040; // @[OneHot.scala 66:30:@2390.4]
  wire [15:0] _T_5081; // @[Mux.scala 31:69:@2408.4]
  wire [15:0] _T_5082; // @[Mux.scala 31:69:@2409.4]
  wire [15:0] _T_5083; // @[Mux.scala 31:69:@2410.4]
  wire [15:0] _T_5084; // @[Mux.scala 31:69:@2411.4]
  wire [15:0] _T_5085; // @[Mux.scala 31:69:@2412.4]
  wire [15:0] _T_5086; // @[Mux.scala 31:69:@2413.4]
  wire [15:0] _T_5087; // @[Mux.scala 31:69:@2414.4]
  wire [15:0] _T_5088; // @[Mux.scala 31:69:@2415.4]
  wire [15:0] _T_5089; // @[Mux.scala 31:69:@2416.4]
  wire [15:0] _T_5090; // @[Mux.scala 31:69:@2417.4]
  wire [15:0] _T_5091; // @[Mux.scala 31:69:@2418.4]
  wire [15:0] _T_5092; // @[Mux.scala 31:69:@2419.4]
  wire [15:0] _T_5093; // @[Mux.scala 31:69:@2420.4]
  wire [15:0] _T_5094; // @[Mux.scala 31:69:@2421.4]
  wire [15:0] _T_5095; // @[Mux.scala 31:69:@2422.4]
  wire [15:0] _T_5096; // @[Mux.scala 31:69:@2423.4]
  wire  _T_5097; // @[OneHot.scala 66:30:@2424.4]
  wire  _T_5098; // @[OneHot.scala 66:30:@2425.4]
  wire  _T_5099; // @[OneHot.scala 66:30:@2426.4]
  wire  _T_5100; // @[OneHot.scala 66:30:@2427.4]
  wire  _T_5101; // @[OneHot.scala 66:30:@2428.4]
  wire  _T_5102; // @[OneHot.scala 66:30:@2429.4]
  wire  _T_5103; // @[OneHot.scala 66:30:@2430.4]
  wire  _T_5104; // @[OneHot.scala 66:30:@2431.4]
  wire  _T_5105; // @[OneHot.scala 66:30:@2432.4]
  wire  _T_5106; // @[OneHot.scala 66:30:@2433.4]
  wire  _T_5107; // @[OneHot.scala 66:30:@2434.4]
  wire  _T_5108; // @[OneHot.scala 66:30:@2435.4]
  wire  _T_5109; // @[OneHot.scala 66:30:@2436.4]
  wire  _T_5110; // @[OneHot.scala 66:30:@2437.4]
  wire  _T_5111; // @[OneHot.scala 66:30:@2438.4]
  wire  _T_5112; // @[OneHot.scala 66:30:@2439.4]
  wire [15:0] _T_5153; // @[Mux.scala 31:69:@2457.4]
  wire [15:0] _T_5154; // @[Mux.scala 31:69:@2458.4]
  wire [15:0] _T_5155; // @[Mux.scala 31:69:@2459.4]
  wire [15:0] _T_5156; // @[Mux.scala 31:69:@2460.4]
  wire [15:0] _T_5157; // @[Mux.scala 31:69:@2461.4]
  wire [15:0] _T_5158; // @[Mux.scala 31:69:@2462.4]
  wire [15:0] _T_5159; // @[Mux.scala 31:69:@2463.4]
  wire [15:0] _T_5160; // @[Mux.scala 31:69:@2464.4]
  wire [15:0] _T_5161; // @[Mux.scala 31:69:@2465.4]
  wire [15:0] _T_5162; // @[Mux.scala 31:69:@2466.4]
  wire [15:0] _T_5163; // @[Mux.scala 31:69:@2467.4]
  wire [15:0] _T_5164; // @[Mux.scala 31:69:@2468.4]
  wire [15:0] _T_5165; // @[Mux.scala 31:69:@2469.4]
  wire [15:0] _T_5166; // @[Mux.scala 31:69:@2470.4]
  wire [15:0] _T_5167; // @[Mux.scala 31:69:@2471.4]
  wire [15:0] _T_5168; // @[Mux.scala 31:69:@2472.4]
  wire  _T_5169; // @[OneHot.scala 66:30:@2473.4]
  wire  _T_5170; // @[OneHot.scala 66:30:@2474.4]
  wire  _T_5171; // @[OneHot.scala 66:30:@2475.4]
  wire  _T_5172; // @[OneHot.scala 66:30:@2476.4]
  wire  _T_5173; // @[OneHot.scala 66:30:@2477.4]
  wire  _T_5174; // @[OneHot.scala 66:30:@2478.4]
  wire  _T_5175; // @[OneHot.scala 66:30:@2479.4]
  wire  _T_5176; // @[OneHot.scala 66:30:@2480.4]
  wire  _T_5177; // @[OneHot.scala 66:30:@2481.4]
  wire  _T_5178; // @[OneHot.scala 66:30:@2482.4]
  wire  _T_5179; // @[OneHot.scala 66:30:@2483.4]
  wire  _T_5180; // @[OneHot.scala 66:30:@2484.4]
  wire  _T_5181; // @[OneHot.scala 66:30:@2485.4]
  wire  _T_5182; // @[OneHot.scala 66:30:@2486.4]
  wire  _T_5183; // @[OneHot.scala 66:30:@2487.4]
  wire  _T_5184; // @[OneHot.scala 66:30:@2488.4]
  wire [15:0] _T_5225; // @[Mux.scala 31:69:@2506.4]
  wire [15:0] _T_5226; // @[Mux.scala 31:69:@2507.4]
  wire [15:0] _T_5227; // @[Mux.scala 31:69:@2508.4]
  wire [15:0] _T_5228; // @[Mux.scala 31:69:@2509.4]
  wire [15:0] _T_5229; // @[Mux.scala 31:69:@2510.4]
  wire [15:0] _T_5230; // @[Mux.scala 31:69:@2511.4]
  wire [15:0] _T_5231; // @[Mux.scala 31:69:@2512.4]
  wire [15:0] _T_5232; // @[Mux.scala 31:69:@2513.4]
  wire [15:0] _T_5233; // @[Mux.scala 31:69:@2514.4]
  wire [15:0] _T_5234; // @[Mux.scala 31:69:@2515.4]
  wire [15:0] _T_5235; // @[Mux.scala 31:69:@2516.4]
  wire [15:0] _T_5236; // @[Mux.scala 31:69:@2517.4]
  wire [15:0] _T_5237; // @[Mux.scala 31:69:@2518.4]
  wire [15:0] _T_5238; // @[Mux.scala 31:69:@2519.4]
  wire [15:0] _T_5239; // @[Mux.scala 31:69:@2520.4]
  wire [15:0] _T_5240; // @[Mux.scala 31:69:@2521.4]
  wire  _T_5241; // @[OneHot.scala 66:30:@2522.4]
  wire  _T_5242; // @[OneHot.scala 66:30:@2523.4]
  wire  _T_5243; // @[OneHot.scala 66:30:@2524.4]
  wire  _T_5244; // @[OneHot.scala 66:30:@2525.4]
  wire  _T_5245; // @[OneHot.scala 66:30:@2526.4]
  wire  _T_5246; // @[OneHot.scala 66:30:@2527.4]
  wire  _T_5247; // @[OneHot.scala 66:30:@2528.4]
  wire  _T_5248; // @[OneHot.scala 66:30:@2529.4]
  wire  _T_5249; // @[OneHot.scala 66:30:@2530.4]
  wire  _T_5250; // @[OneHot.scala 66:30:@2531.4]
  wire  _T_5251; // @[OneHot.scala 66:30:@2532.4]
  wire  _T_5252; // @[OneHot.scala 66:30:@2533.4]
  wire  _T_5253; // @[OneHot.scala 66:30:@2534.4]
  wire  _T_5254; // @[OneHot.scala 66:30:@2535.4]
  wire  _T_5255; // @[OneHot.scala 66:30:@2536.4]
  wire  _T_5256; // @[OneHot.scala 66:30:@2537.4]
  wire [15:0] _T_5297; // @[Mux.scala 31:69:@2555.4]
  wire [15:0] _T_5298; // @[Mux.scala 31:69:@2556.4]
  wire [15:0] _T_5299; // @[Mux.scala 31:69:@2557.4]
  wire [15:0] _T_5300; // @[Mux.scala 31:69:@2558.4]
  wire [15:0] _T_5301; // @[Mux.scala 31:69:@2559.4]
  wire [15:0] _T_5302; // @[Mux.scala 31:69:@2560.4]
  wire [15:0] _T_5303; // @[Mux.scala 31:69:@2561.4]
  wire [15:0] _T_5304; // @[Mux.scala 31:69:@2562.4]
  wire [15:0] _T_5305; // @[Mux.scala 31:69:@2563.4]
  wire [15:0] _T_5306; // @[Mux.scala 31:69:@2564.4]
  wire [15:0] _T_5307; // @[Mux.scala 31:69:@2565.4]
  wire [15:0] _T_5308; // @[Mux.scala 31:69:@2566.4]
  wire [15:0] _T_5309; // @[Mux.scala 31:69:@2567.4]
  wire [15:0] _T_5310; // @[Mux.scala 31:69:@2568.4]
  wire [15:0] _T_5311; // @[Mux.scala 31:69:@2569.4]
  wire [15:0] _T_5312; // @[Mux.scala 31:69:@2570.4]
  wire  _T_5313; // @[OneHot.scala 66:30:@2571.4]
  wire  _T_5314; // @[OneHot.scala 66:30:@2572.4]
  wire  _T_5315; // @[OneHot.scala 66:30:@2573.4]
  wire  _T_5316; // @[OneHot.scala 66:30:@2574.4]
  wire  _T_5317; // @[OneHot.scala 66:30:@2575.4]
  wire  _T_5318; // @[OneHot.scala 66:30:@2576.4]
  wire  _T_5319; // @[OneHot.scala 66:30:@2577.4]
  wire  _T_5320; // @[OneHot.scala 66:30:@2578.4]
  wire  _T_5321; // @[OneHot.scala 66:30:@2579.4]
  wire  _T_5322; // @[OneHot.scala 66:30:@2580.4]
  wire  _T_5323; // @[OneHot.scala 66:30:@2581.4]
  wire  _T_5324; // @[OneHot.scala 66:30:@2582.4]
  wire  _T_5325; // @[OneHot.scala 66:30:@2583.4]
  wire  _T_5326; // @[OneHot.scala 66:30:@2584.4]
  wire  _T_5327; // @[OneHot.scala 66:30:@2585.4]
  wire  _T_5328; // @[OneHot.scala 66:30:@2586.4]
  wire [15:0] _T_5369; // @[Mux.scala 31:69:@2604.4]
  wire [15:0] _T_5370; // @[Mux.scala 31:69:@2605.4]
  wire [15:0] _T_5371; // @[Mux.scala 31:69:@2606.4]
  wire [15:0] _T_5372; // @[Mux.scala 31:69:@2607.4]
  wire [15:0] _T_5373; // @[Mux.scala 31:69:@2608.4]
  wire [15:0] _T_5374; // @[Mux.scala 31:69:@2609.4]
  wire [15:0] _T_5375; // @[Mux.scala 31:69:@2610.4]
  wire [15:0] _T_5376; // @[Mux.scala 31:69:@2611.4]
  wire [15:0] _T_5377; // @[Mux.scala 31:69:@2612.4]
  wire [15:0] _T_5378; // @[Mux.scala 31:69:@2613.4]
  wire [15:0] _T_5379; // @[Mux.scala 31:69:@2614.4]
  wire [15:0] _T_5380; // @[Mux.scala 31:69:@2615.4]
  wire [15:0] _T_5381; // @[Mux.scala 31:69:@2616.4]
  wire [15:0] _T_5382; // @[Mux.scala 31:69:@2617.4]
  wire [15:0] _T_5383; // @[Mux.scala 31:69:@2618.4]
  wire [15:0] _T_5384; // @[Mux.scala 31:69:@2619.4]
  wire  _T_5385; // @[OneHot.scala 66:30:@2620.4]
  wire  _T_5386; // @[OneHot.scala 66:30:@2621.4]
  wire  _T_5387; // @[OneHot.scala 66:30:@2622.4]
  wire  _T_5388; // @[OneHot.scala 66:30:@2623.4]
  wire  _T_5389; // @[OneHot.scala 66:30:@2624.4]
  wire  _T_5390; // @[OneHot.scala 66:30:@2625.4]
  wire  _T_5391; // @[OneHot.scala 66:30:@2626.4]
  wire  _T_5392; // @[OneHot.scala 66:30:@2627.4]
  wire  _T_5393; // @[OneHot.scala 66:30:@2628.4]
  wire  _T_5394; // @[OneHot.scala 66:30:@2629.4]
  wire  _T_5395; // @[OneHot.scala 66:30:@2630.4]
  wire  _T_5396; // @[OneHot.scala 66:30:@2631.4]
  wire  _T_5397; // @[OneHot.scala 66:30:@2632.4]
  wire  _T_5398; // @[OneHot.scala 66:30:@2633.4]
  wire  _T_5399; // @[OneHot.scala 66:30:@2634.4]
  wire  _T_5400; // @[OneHot.scala 66:30:@2635.4]
  wire [15:0] _T_5441; // @[Mux.scala 31:69:@2653.4]
  wire [15:0] _T_5442; // @[Mux.scala 31:69:@2654.4]
  wire [15:0] _T_5443; // @[Mux.scala 31:69:@2655.4]
  wire [15:0] _T_5444; // @[Mux.scala 31:69:@2656.4]
  wire [15:0] _T_5445; // @[Mux.scala 31:69:@2657.4]
  wire [15:0] _T_5446; // @[Mux.scala 31:69:@2658.4]
  wire [15:0] _T_5447; // @[Mux.scala 31:69:@2659.4]
  wire [15:0] _T_5448; // @[Mux.scala 31:69:@2660.4]
  wire [15:0] _T_5449; // @[Mux.scala 31:69:@2661.4]
  wire [15:0] _T_5450; // @[Mux.scala 31:69:@2662.4]
  wire [15:0] _T_5451; // @[Mux.scala 31:69:@2663.4]
  wire [15:0] _T_5452; // @[Mux.scala 31:69:@2664.4]
  wire [15:0] _T_5453; // @[Mux.scala 31:69:@2665.4]
  wire [15:0] _T_5454; // @[Mux.scala 31:69:@2666.4]
  wire [15:0] _T_5455; // @[Mux.scala 31:69:@2667.4]
  wire [15:0] _T_5456; // @[Mux.scala 31:69:@2668.4]
  wire  _T_5457; // @[OneHot.scala 66:30:@2669.4]
  wire  _T_5458; // @[OneHot.scala 66:30:@2670.4]
  wire  _T_5459; // @[OneHot.scala 66:30:@2671.4]
  wire  _T_5460; // @[OneHot.scala 66:30:@2672.4]
  wire  _T_5461; // @[OneHot.scala 66:30:@2673.4]
  wire  _T_5462; // @[OneHot.scala 66:30:@2674.4]
  wire  _T_5463; // @[OneHot.scala 66:30:@2675.4]
  wire  _T_5464; // @[OneHot.scala 66:30:@2676.4]
  wire  _T_5465; // @[OneHot.scala 66:30:@2677.4]
  wire  _T_5466; // @[OneHot.scala 66:30:@2678.4]
  wire  _T_5467; // @[OneHot.scala 66:30:@2679.4]
  wire  _T_5468; // @[OneHot.scala 66:30:@2680.4]
  wire  _T_5469; // @[OneHot.scala 66:30:@2681.4]
  wire  _T_5470; // @[OneHot.scala 66:30:@2682.4]
  wire  _T_5471; // @[OneHot.scala 66:30:@2683.4]
  wire  _T_5472; // @[OneHot.scala 66:30:@2684.4]
  wire [15:0] _T_5513; // @[Mux.scala 31:69:@2702.4]
  wire [15:0] _T_5514; // @[Mux.scala 31:69:@2703.4]
  wire [15:0] _T_5515; // @[Mux.scala 31:69:@2704.4]
  wire [15:0] _T_5516; // @[Mux.scala 31:69:@2705.4]
  wire [15:0] _T_5517; // @[Mux.scala 31:69:@2706.4]
  wire [15:0] _T_5518; // @[Mux.scala 31:69:@2707.4]
  wire [15:0] _T_5519; // @[Mux.scala 31:69:@2708.4]
  wire [15:0] _T_5520; // @[Mux.scala 31:69:@2709.4]
  wire [15:0] _T_5521; // @[Mux.scala 31:69:@2710.4]
  wire [15:0] _T_5522; // @[Mux.scala 31:69:@2711.4]
  wire [15:0] _T_5523; // @[Mux.scala 31:69:@2712.4]
  wire [15:0] _T_5524; // @[Mux.scala 31:69:@2713.4]
  wire [15:0] _T_5525; // @[Mux.scala 31:69:@2714.4]
  wire [15:0] _T_5526; // @[Mux.scala 31:69:@2715.4]
  wire [15:0] _T_5527; // @[Mux.scala 31:69:@2716.4]
  wire [15:0] _T_5528; // @[Mux.scala 31:69:@2717.4]
  wire  _T_5529; // @[OneHot.scala 66:30:@2718.4]
  wire  _T_5530; // @[OneHot.scala 66:30:@2719.4]
  wire  _T_5531; // @[OneHot.scala 66:30:@2720.4]
  wire  _T_5532; // @[OneHot.scala 66:30:@2721.4]
  wire  _T_5533; // @[OneHot.scala 66:30:@2722.4]
  wire  _T_5534; // @[OneHot.scala 66:30:@2723.4]
  wire  _T_5535; // @[OneHot.scala 66:30:@2724.4]
  wire  _T_5536; // @[OneHot.scala 66:30:@2725.4]
  wire  _T_5537; // @[OneHot.scala 66:30:@2726.4]
  wire  _T_5538; // @[OneHot.scala 66:30:@2727.4]
  wire  _T_5539; // @[OneHot.scala 66:30:@2728.4]
  wire  _T_5540; // @[OneHot.scala 66:30:@2729.4]
  wire  _T_5541; // @[OneHot.scala 66:30:@2730.4]
  wire  _T_5542; // @[OneHot.scala 66:30:@2731.4]
  wire  _T_5543; // @[OneHot.scala 66:30:@2732.4]
  wire  _T_5544; // @[OneHot.scala 66:30:@2733.4]
  wire [15:0] _T_5585; // @[Mux.scala 31:69:@2751.4]
  wire [15:0] _T_5586; // @[Mux.scala 31:69:@2752.4]
  wire [15:0] _T_5587; // @[Mux.scala 31:69:@2753.4]
  wire [15:0] _T_5588; // @[Mux.scala 31:69:@2754.4]
  wire [15:0] _T_5589; // @[Mux.scala 31:69:@2755.4]
  wire [15:0] _T_5590; // @[Mux.scala 31:69:@2756.4]
  wire [15:0] _T_5591; // @[Mux.scala 31:69:@2757.4]
  wire [15:0] _T_5592; // @[Mux.scala 31:69:@2758.4]
  wire [15:0] _T_5593; // @[Mux.scala 31:69:@2759.4]
  wire [15:0] _T_5594; // @[Mux.scala 31:69:@2760.4]
  wire [15:0] _T_5595; // @[Mux.scala 31:69:@2761.4]
  wire [15:0] _T_5596; // @[Mux.scala 31:69:@2762.4]
  wire [15:0] _T_5597; // @[Mux.scala 31:69:@2763.4]
  wire [15:0] _T_5598; // @[Mux.scala 31:69:@2764.4]
  wire [15:0] _T_5599; // @[Mux.scala 31:69:@2765.4]
  wire [15:0] _T_5600; // @[Mux.scala 31:69:@2766.4]
  wire  _T_5601; // @[OneHot.scala 66:30:@2767.4]
  wire  _T_5602; // @[OneHot.scala 66:30:@2768.4]
  wire  _T_5603; // @[OneHot.scala 66:30:@2769.4]
  wire  _T_5604; // @[OneHot.scala 66:30:@2770.4]
  wire  _T_5605; // @[OneHot.scala 66:30:@2771.4]
  wire  _T_5606; // @[OneHot.scala 66:30:@2772.4]
  wire  _T_5607; // @[OneHot.scala 66:30:@2773.4]
  wire  _T_5608; // @[OneHot.scala 66:30:@2774.4]
  wire  _T_5609; // @[OneHot.scala 66:30:@2775.4]
  wire  _T_5610; // @[OneHot.scala 66:30:@2776.4]
  wire  _T_5611; // @[OneHot.scala 66:30:@2777.4]
  wire  _T_5612; // @[OneHot.scala 66:30:@2778.4]
  wire  _T_5613; // @[OneHot.scala 66:30:@2779.4]
  wire  _T_5614; // @[OneHot.scala 66:30:@2780.4]
  wire  _T_5615; // @[OneHot.scala 66:30:@2781.4]
  wire  _T_5616; // @[OneHot.scala 66:30:@2782.4]
  wire [15:0] _T_5657; // @[Mux.scala 31:69:@2800.4]
  wire [15:0] _T_5658; // @[Mux.scala 31:69:@2801.4]
  wire [15:0] _T_5659; // @[Mux.scala 31:69:@2802.4]
  wire [15:0] _T_5660; // @[Mux.scala 31:69:@2803.4]
  wire [15:0] _T_5661; // @[Mux.scala 31:69:@2804.4]
  wire [15:0] _T_5662; // @[Mux.scala 31:69:@2805.4]
  wire [15:0] _T_5663; // @[Mux.scala 31:69:@2806.4]
  wire [15:0] _T_5664; // @[Mux.scala 31:69:@2807.4]
  wire [15:0] _T_5665; // @[Mux.scala 31:69:@2808.4]
  wire [15:0] _T_5666; // @[Mux.scala 31:69:@2809.4]
  wire [15:0] _T_5667; // @[Mux.scala 31:69:@2810.4]
  wire [15:0] _T_5668; // @[Mux.scala 31:69:@2811.4]
  wire [15:0] _T_5669; // @[Mux.scala 31:69:@2812.4]
  wire [15:0] _T_5670; // @[Mux.scala 31:69:@2813.4]
  wire [15:0] _T_5671; // @[Mux.scala 31:69:@2814.4]
  wire [15:0] _T_5672; // @[Mux.scala 31:69:@2815.4]
  wire  _T_5673; // @[OneHot.scala 66:30:@2816.4]
  wire  _T_5674; // @[OneHot.scala 66:30:@2817.4]
  wire  _T_5675; // @[OneHot.scala 66:30:@2818.4]
  wire  _T_5676; // @[OneHot.scala 66:30:@2819.4]
  wire  _T_5677; // @[OneHot.scala 66:30:@2820.4]
  wire  _T_5678; // @[OneHot.scala 66:30:@2821.4]
  wire  _T_5679; // @[OneHot.scala 66:30:@2822.4]
  wire  _T_5680; // @[OneHot.scala 66:30:@2823.4]
  wire  _T_5681; // @[OneHot.scala 66:30:@2824.4]
  wire  _T_5682; // @[OneHot.scala 66:30:@2825.4]
  wire  _T_5683; // @[OneHot.scala 66:30:@2826.4]
  wire  _T_5684; // @[OneHot.scala 66:30:@2827.4]
  wire  _T_5685; // @[OneHot.scala 66:30:@2828.4]
  wire  _T_5686; // @[OneHot.scala 66:30:@2829.4]
  wire  _T_5687; // @[OneHot.scala 66:30:@2830.4]
  wire  _T_5688; // @[OneHot.scala 66:30:@2831.4]
  wire [7:0] _T_5753; // @[Mux.scala 19:72:@2855.4]
  wire [15:0] _T_5761; // @[Mux.scala 19:72:@2863.4]
  wire [15:0] _T_5763; // @[Mux.scala 19:72:@2864.4]
  wire [7:0] _T_5770; // @[Mux.scala 19:72:@2871.4]
  wire [15:0] _T_5778; // @[Mux.scala 19:72:@2879.4]
  wire [15:0] _T_5780; // @[Mux.scala 19:72:@2880.4]
  wire [7:0] _T_5787; // @[Mux.scala 19:72:@2887.4]
  wire [15:0] _T_5795; // @[Mux.scala 19:72:@2895.4]
  wire [15:0] _T_5797; // @[Mux.scala 19:72:@2896.4]
  wire [7:0] _T_5804; // @[Mux.scala 19:72:@2903.4]
  wire [15:0] _T_5812; // @[Mux.scala 19:72:@2911.4]
  wire [15:0] _T_5814; // @[Mux.scala 19:72:@2912.4]
  wire [7:0] _T_5821; // @[Mux.scala 19:72:@2919.4]
  wire [15:0] _T_5829; // @[Mux.scala 19:72:@2927.4]
  wire [15:0] _T_5831; // @[Mux.scala 19:72:@2928.4]
  wire [7:0] _T_5838; // @[Mux.scala 19:72:@2935.4]
  wire [15:0] _T_5846; // @[Mux.scala 19:72:@2943.4]
  wire [15:0] _T_5848; // @[Mux.scala 19:72:@2944.4]
  wire [7:0] _T_5855; // @[Mux.scala 19:72:@2951.4]
  wire [15:0] _T_5863; // @[Mux.scala 19:72:@2959.4]
  wire [15:0] _T_5865; // @[Mux.scala 19:72:@2960.4]
  wire [7:0] _T_5872; // @[Mux.scala 19:72:@2967.4]
  wire [15:0] _T_5880; // @[Mux.scala 19:72:@2975.4]
  wire [15:0] _T_5882; // @[Mux.scala 19:72:@2976.4]
  wire [7:0] _T_5889; // @[Mux.scala 19:72:@2983.4]
  wire [15:0] _T_5897; // @[Mux.scala 19:72:@2991.4]
  wire [15:0] _T_5899; // @[Mux.scala 19:72:@2992.4]
  wire [7:0] _T_5906; // @[Mux.scala 19:72:@2999.4]
  wire [15:0] _T_5914; // @[Mux.scala 19:72:@3007.4]
  wire [15:0] _T_5916; // @[Mux.scala 19:72:@3008.4]
  wire [7:0] _T_5923; // @[Mux.scala 19:72:@3015.4]
  wire [15:0] _T_5931; // @[Mux.scala 19:72:@3023.4]
  wire [15:0] _T_5933; // @[Mux.scala 19:72:@3024.4]
  wire [7:0] _T_5940; // @[Mux.scala 19:72:@3031.4]
  wire [15:0] _T_5948; // @[Mux.scala 19:72:@3039.4]
  wire [15:0] _T_5950; // @[Mux.scala 19:72:@3040.4]
  wire [7:0] _T_5957; // @[Mux.scala 19:72:@3047.4]
  wire [15:0] _T_5965; // @[Mux.scala 19:72:@3055.4]
  wire [15:0] _T_5967; // @[Mux.scala 19:72:@3056.4]
  wire [7:0] _T_5974; // @[Mux.scala 19:72:@3063.4]
  wire [15:0] _T_5982; // @[Mux.scala 19:72:@3071.4]
  wire [15:0] _T_5984; // @[Mux.scala 19:72:@3072.4]
  wire [7:0] _T_5991; // @[Mux.scala 19:72:@3079.4]
  wire [15:0] _T_5999; // @[Mux.scala 19:72:@3087.4]
  wire [15:0] _T_6001; // @[Mux.scala 19:72:@3088.4]
  wire [7:0] _T_6008; // @[Mux.scala 19:72:@3095.4]
  wire [15:0] _T_6016; // @[Mux.scala 19:72:@3103.4]
  wire [15:0] _T_6018; // @[Mux.scala 19:72:@3104.4]
  wire [15:0] _T_6019; // @[Mux.scala 19:72:@3105.4]
  wire [15:0] _T_6020; // @[Mux.scala 19:72:@3106.4]
  wire [15:0] _T_6021; // @[Mux.scala 19:72:@3107.4]
  wire [15:0] _T_6022; // @[Mux.scala 19:72:@3108.4]
  wire [15:0] _T_6023; // @[Mux.scala 19:72:@3109.4]
  wire [15:0] _T_6024; // @[Mux.scala 19:72:@3110.4]
  wire [15:0] _T_6025; // @[Mux.scala 19:72:@3111.4]
  wire [15:0] _T_6026; // @[Mux.scala 19:72:@3112.4]
  wire [15:0] _T_6027; // @[Mux.scala 19:72:@3113.4]
  wire [15:0] _T_6028; // @[Mux.scala 19:72:@3114.4]
  wire [15:0] _T_6029; // @[Mux.scala 19:72:@3115.4]
  wire [15:0] _T_6030; // @[Mux.scala 19:72:@3116.4]
  wire [15:0] _T_6031; // @[Mux.scala 19:72:@3117.4]
  wire [15:0] _T_6032; // @[Mux.scala 19:72:@3118.4]
  wire [15:0] _T_6033; // @[Mux.scala 19:72:@3119.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@3123.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@3125.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@3127.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@3129.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@3131.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@3133.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@3135.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@3137.4]
  wire  inputAddrPriorityPorts_0_8; // @[Mux.scala 19:72:@3139.4]
  wire  inputAddrPriorityPorts_0_9; // @[Mux.scala 19:72:@3141.4]
  wire  inputAddrPriorityPorts_0_10; // @[Mux.scala 19:72:@3143.4]
  wire  inputAddrPriorityPorts_0_11; // @[Mux.scala 19:72:@3145.4]
  wire  inputAddrPriorityPorts_0_12; // @[Mux.scala 19:72:@3147.4]
  wire  inputAddrPriorityPorts_0_13; // @[Mux.scala 19:72:@3149.4]
  wire  inputAddrPriorityPorts_0_14; // @[Mux.scala 19:72:@3151.4]
  wire  inputAddrPriorityPorts_0_15; // @[Mux.scala 19:72:@3153.4]
  wire [15:0] _T_6235; // @[Mux.scala 31:69:@3207.4]
  wire [15:0] _T_6236; // @[Mux.scala 31:69:@3208.4]
  wire [15:0] _T_6237; // @[Mux.scala 31:69:@3209.4]
  wire [15:0] _T_6238; // @[Mux.scala 31:69:@3210.4]
  wire [15:0] _T_6239; // @[Mux.scala 31:69:@3211.4]
  wire [15:0] _T_6240; // @[Mux.scala 31:69:@3212.4]
  wire [15:0] _T_6241; // @[Mux.scala 31:69:@3213.4]
  wire [15:0] _T_6242; // @[Mux.scala 31:69:@3214.4]
  wire [15:0] _T_6243; // @[Mux.scala 31:69:@3215.4]
  wire [15:0] _T_6244; // @[Mux.scala 31:69:@3216.4]
  wire [15:0] _T_6245; // @[Mux.scala 31:69:@3217.4]
  wire [15:0] _T_6246; // @[Mux.scala 31:69:@3218.4]
  wire [15:0] _T_6247; // @[Mux.scala 31:69:@3219.4]
  wire [15:0] _T_6248; // @[Mux.scala 31:69:@3220.4]
  wire [15:0] _T_6249; // @[Mux.scala 31:69:@3221.4]
  wire [15:0] _T_6250; // @[Mux.scala 31:69:@3222.4]
  wire  _T_6251; // @[OneHot.scala 66:30:@3223.4]
  wire  _T_6252; // @[OneHot.scala 66:30:@3224.4]
  wire  _T_6253; // @[OneHot.scala 66:30:@3225.4]
  wire  _T_6254; // @[OneHot.scala 66:30:@3226.4]
  wire  _T_6255; // @[OneHot.scala 66:30:@3227.4]
  wire  _T_6256; // @[OneHot.scala 66:30:@3228.4]
  wire  _T_6257; // @[OneHot.scala 66:30:@3229.4]
  wire  _T_6258; // @[OneHot.scala 66:30:@3230.4]
  wire  _T_6259; // @[OneHot.scala 66:30:@3231.4]
  wire  _T_6260; // @[OneHot.scala 66:30:@3232.4]
  wire  _T_6261; // @[OneHot.scala 66:30:@3233.4]
  wire  _T_6262; // @[OneHot.scala 66:30:@3234.4]
  wire  _T_6263; // @[OneHot.scala 66:30:@3235.4]
  wire  _T_6264; // @[OneHot.scala 66:30:@3236.4]
  wire  _T_6265; // @[OneHot.scala 66:30:@3237.4]
  wire  _T_6266; // @[OneHot.scala 66:30:@3238.4]
  wire [15:0] _T_6307; // @[Mux.scala 31:69:@3256.4]
  wire [15:0] _T_6308; // @[Mux.scala 31:69:@3257.4]
  wire [15:0] _T_6309; // @[Mux.scala 31:69:@3258.4]
  wire [15:0] _T_6310; // @[Mux.scala 31:69:@3259.4]
  wire [15:0] _T_6311; // @[Mux.scala 31:69:@3260.4]
  wire [15:0] _T_6312; // @[Mux.scala 31:69:@3261.4]
  wire [15:0] _T_6313; // @[Mux.scala 31:69:@3262.4]
  wire [15:0] _T_6314; // @[Mux.scala 31:69:@3263.4]
  wire [15:0] _T_6315; // @[Mux.scala 31:69:@3264.4]
  wire [15:0] _T_6316; // @[Mux.scala 31:69:@3265.4]
  wire [15:0] _T_6317; // @[Mux.scala 31:69:@3266.4]
  wire [15:0] _T_6318; // @[Mux.scala 31:69:@3267.4]
  wire [15:0] _T_6319; // @[Mux.scala 31:69:@3268.4]
  wire [15:0] _T_6320; // @[Mux.scala 31:69:@3269.4]
  wire [15:0] _T_6321; // @[Mux.scala 31:69:@3270.4]
  wire [15:0] _T_6322; // @[Mux.scala 31:69:@3271.4]
  wire  _T_6323; // @[OneHot.scala 66:30:@3272.4]
  wire  _T_6324; // @[OneHot.scala 66:30:@3273.4]
  wire  _T_6325; // @[OneHot.scala 66:30:@3274.4]
  wire  _T_6326; // @[OneHot.scala 66:30:@3275.4]
  wire  _T_6327; // @[OneHot.scala 66:30:@3276.4]
  wire  _T_6328; // @[OneHot.scala 66:30:@3277.4]
  wire  _T_6329; // @[OneHot.scala 66:30:@3278.4]
  wire  _T_6330; // @[OneHot.scala 66:30:@3279.4]
  wire  _T_6331; // @[OneHot.scala 66:30:@3280.4]
  wire  _T_6332; // @[OneHot.scala 66:30:@3281.4]
  wire  _T_6333; // @[OneHot.scala 66:30:@3282.4]
  wire  _T_6334; // @[OneHot.scala 66:30:@3283.4]
  wire  _T_6335; // @[OneHot.scala 66:30:@3284.4]
  wire  _T_6336; // @[OneHot.scala 66:30:@3285.4]
  wire  _T_6337; // @[OneHot.scala 66:30:@3286.4]
  wire  _T_6338; // @[OneHot.scala 66:30:@3287.4]
  wire [15:0] _T_6379; // @[Mux.scala 31:69:@3305.4]
  wire [15:0] _T_6380; // @[Mux.scala 31:69:@3306.4]
  wire [15:0] _T_6381; // @[Mux.scala 31:69:@3307.4]
  wire [15:0] _T_6382; // @[Mux.scala 31:69:@3308.4]
  wire [15:0] _T_6383; // @[Mux.scala 31:69:@3309.4]
  wire [15:0] _T_6384; // @[Mux.scala 31:69:@3310.4]
  wire [15:0] _T_6385; // @[Mux.scala 31:69:@3311.4]
  wire [15:0] _T_6386; // @[Mux.scala 31:69:@3312.4]
  wire [15:0] _T_6387; // @[Mux.scala 31:69:@3313.4]
  wire [15:0] _T_6388; // @[Mux.scala 31:69:@3314.4]
  wire [15:0] _T_6389; // @[Mux.scala 31:69:@3315.4]
  wire [15:0] _T_6390; // @[Mux.scala 31:69:@3316.4]
  wire [15:0] _T_6391; // @[Mux.scala 31:69:@3317.4]
  wire [15:0] _T_6392; // @[Mux.scala 31:69:@3318.4]
  wire [15:0] _T_6393; // @[Mux.scala 31:69:@3319.4]
  wire [15:0] _T_6394; // @[Mux.scala 31:69:@3320.4]
  wire  _T_6395; // @[OneHot.scala 66:30:@3321.4]
  wire  _T_6396; // @[OneHot.scala 66:30:@3322.4]
  wire  _T_6397; // @[OneHot.scala 66:30:@3323.4]
  wire  _T_6398; // @[OneHot.scala 66:30:@3324.4]
  wire  _T_6399; // @[OneHot.scala 66:30:@3325.4]
  wire  _T_6400; // @[OneHot.scala 66:30:@3326.4]
  wire  _T_6401; // @[OneHot.scala 66:30:@3327.4]
  wire  _T_6402; // @[OneHot.scala 66:30:@3328.4]
  wire  _T_6403; // @[OneHot.scala 66:30:@3329.4]
  wire  _T_6404; // @[OneHot.scala 66:30:@3330.4]
  wire  _T_6405; // @[OneHot.scala 66:30:@3331.4]
  wire  _T_6406; // @[OneHot.scala 66:30:@3332.4]
  wire  _T_6407; // @[OneHot.scala 66:30:@3333.4]
  wire  _T_6408; // @[OneHot.scala 66:30:@3334.4]
  wire  _T_6409; // @[OneHot.scala 66:30:@3335.4]
  wire  _T_6410; // @[OneHot.scala 66:30:@3336.4]
  wire [15:0] _T_6451; // @[Mux.scala 31:69:@3354.4]
  wire [15:0] _T_6452; // @[Mux.scala 31:69:@3355.4]
  wire [15:0] _T_6453; // @[Mux.scala 31:69:@3356.4]
  wire [15:0] _T_6454; // @[Mux.scala 31:69:@3357.4]
  wire [15:0] _T_6455; // @[Mux.scala 31:69:@3358.4]
  wire [15:0] _T_6456; // @[Mux.scala 31:69:@3359.4]
  wire [15:0] _T_6457; // @[Mux.scala 31:69:@3360.4]
  wire [15:0] _T_6458; // @[Mux.scala 31:69:@3361.4]
  wire [15:0] _T_6459; // @[Mux.scala 31:69:@3362.4]
  wire [15:0] _T_6460; // @[Mux.scala 31:69:@3363.4]
  wire [15:0] _T_6461; // @[Mux.scala 31:69:@3364.4]
  wire [15:0] _T_6462; // @[Mux.scala 31:69:@3365.4]
  wire [15:0] _T_6463; // @[Mux.scala 31:69:@3366.4]
  wire [15:0] _T_6464; // @[Mux.scala 31:69:@3367.4]
  wire [15:0] _T_6465; // @[Mux.scala 31:69:@3368.4]
  wire [15:0] _T_6466; // @[Mux.scala 31:69:@3369.4]
  wire  _T_6467; // @[OneHot.scala 66:30:@3370.4]
  wire  _T_6468; // @[OneHot.scala 66:30:@3371.4]
  wire  _T_6469; // @[OneHot.scala 66:30:@3372.4]
  wire  _T_6470; // @[OneHot.scala 66:30:@3373.4]
  wire  _T_6471; // @[OneHot.scala 66:30:@3374.4]
  wire  _T_6472; // @[OneHot.scala 66:30:@3375.4]
  wire  _T_6473; // @[OneHot.scala 66:30:@3376.4]
  wire  _T_6474; // @[OneHot.scala 66:30:@3377.4]
  wire  _T_6475; // @[OneHot.scala 66:30:@3378.4]
  wire  _T_6476; // @[OneHot.scala 66:30:@3379.4]
  wire  _T_6477; // @[OneHot.scala 66:30:@3380.4]
  wire  _T_6478; // @[OneHot.scala 66:30:@3381.4]
  wire  _T_6479; // @[OneHot.scala 66:30:@3382.4]
  wire  _T_6480; // @[OneHot.scala 66:30:@3383.4]
  wire  _T_6481; // @[OneHot.scala 66:30:@3384.4]
  wire  _T_6482; // @[OneHot.scala 66:30:@3385.4]
  wire [15:0] _T_6523; // @[Mux.scala 31:69:@3403.4]
  wire [15:0] _T_6524; // @[Mux.scala 31:69:@3404.4]
  wire [15:0] _T_6525; // @[Mux.scala 31:69:@3405.4]
  wire [15:0] _T_6526; // @[Mux.scala 31:69:@3406.4]
  wire [15:0] _T_6527; // @[Mux.scala 31:69:@3407.4]
  wire [15:0] _T_6528; // @[Mux.scala 31:69:@3408.4]
  wire [15:0] _T_6529; // @[Mux.scala 31:69:@3409.4]
  wire [15:0] _T_6530; // @[Mux.scala 31:69:@3410.4]
  wire [15:0] _T_6531; // @[Mux.scala 31:69:@3411.4]
  wire [15:0] _T_6532; // @[Mux.scala 31:69:@3412.4]
  wire [15:0] _T_6533; // @[Mux.scala 31:69:@3413.4]
  wire [15:0] _T_6534; // @[Mux.scala 31:69:@3414.4]
  wire [15:0] _T_6535; // @[Mux.scala 31:69:@3415.4]
  wire [15:0] _T_6536; // @[Mux.scala 31:69:@3416.4]
  wire [15:0] _T_6537; // @[Mux.scala 31:69:@3417.4]
  wire [15:0] _T_6538; // @[Mux.scala 31:69:@3418.4]
  wire  _T_6539; // @[OneHot.scala 66:30:@3419.4]
  wire  _T_6540; // @[OneHot.scala 66:30:@3420.4]
  wire  _T_6541; // @[OneHot.scala 66:30:@3421.4]
  wire  _T_6542; // @[OneHot.scala 66:30:@3422.4]
  wire  _T_6543; // @[OneHot.scala 66:30:@3423.4]
  wire  _T_6544; // @[OneHot.scala 66:30:@3424.4]
  wire  _T_6545; // @[OneHot.scala 66:30:@3425.4]
  wire  _T_6546; // @[OneHot.scala 66:30:@3426.4]
  wire  _T_6547; // @[OneHot.scala 66:30:@3427.4]
  wire  _T_6548; // @[OneHot.scala 66:30:@3428.4]
  wire  _T_6549; // @[OneHot.scala 66:30:@3429.4]
  wire  _T_6550; // @[OneHot.scala 66:30:@3430.4]
  wire  _T_6551; // @[OneHot.scala 66:30:@3431.4]
  wire  _T_6552; // @[OneHot.scala 66:30:@3432.4]
  wire  _T_6553; // @[OneHot.scala 66:30:@3433.4]
  wire  _T_6554; // @[OneHot.scala 66:30:@3434.4]
  wire [15:0] _T_6595; // @[Mux.scala 31:69:@3452.4]
  wire [15:0] _T_6596; // @[Mux.scala 31:69:@3453.4]
  wire [15:0] _T_6597; // @[Mux.scala 31:69:@3454.4]
  wire [15:0] _T_6598; // @[Mux.scala 31:69:@3455.4]
  wire [15:0] _T_6599; // @[Mux.scala 31:69:@3456.4]
  wire [15:0] _T_6600; // @[Mux.scala 31:69:@3457.4]
  wire [15:0] _T_6601; // @[Mux.scala 31:69:@3458.4]
  wire [15:0] _T_6602; // @[Mux.scala 31:69:@3459.4]
  wire [15:0] _T_6603; // @[Mux.scala 31:69:@3460.4]
  wire [15:0] _T_6604; // @[Mux.scala 31:69:@3461.4]
  wire [15:0] _T_6605; // @[Mux.scala 31:69:@3462.4]
  wire [15:0] _T_6606; // @[Mux.scala 31:69:@3463.4]
  wire [15:0] _T_6607; // @[Mux.scala 31:69:@3464.4]
  wire [15:0] _T_6608; // @[Mux.scala 31:69:@3465.4]
  wire [15:0] _T_6609; // @[Mux.scala 31:69:@3466.4]
  wire [15:0] _T_6610; // @[Mux.scala 31:69:@3467.4]
  wire  _T_6611; // @[OneHot.scala 66:30:@3468.4]
  wire  _T_6612; // @[OneHot.scala 66:30:@3469.4]
  wire  _T_6613; // @[OneHot.scala 66:30:@3470.4]
  wire  _T_6614; // @[OneHot.scala 66:30:@3471.4]
  wire  _T_6615; // @[OneHot.scala 66:30:@3472.4]
  wire  _T_6616; // @[OneHot.scala 66:30:@3473.4]
  wire  _T_6617; // @[OneHot.scala 66:30:@3474.4]
  wire  _T_6618; // @[OneHot.scala 66:30:@3475.4]
  wire  _T_6619; // @[OneHot.scala 66:30:@3476.4]
  wire  _T_6620; // @[OneHot.scala 66:30:@3477.4]
  wire  _T_6621; // @[OneHot.scala 66:30:@3478.4]
  wire  _T_6622; // @[OneHot.scala 66:30:@3479.4]
  wire  _T_6623; // @[OneHot.scala 66:30:@3480.4]
  wire  _T_6624; // @[OneHot.scala 66:30:@3481.4]
  wire  _T_6625; // @[OneHot.scala 66:30:@3482.4]
  wire  _T_6626; // @[OneHot.scala 66:30:@3483.4]
  wire [15:0] _T_6667; // @[Mux.scala 31:69:@3501.4]
  wire [15:0] _T_6668; // @[Mux.scala 31:69:@3502.4]
  wire [15:0] _T_6669; // @[Mux.scala 31:69:@3503.4]
  wire [15:0] _T_6670; // @[Mux.scala 31:69:@3504.4]
  wire [15:0] _T_6671; // @[Mux.scala 31:69:@3505.4]
  wire [15:0] _T_6672; // @[Mux.scala 31:69:@3506.4]
  wire [15:0] _T_6673; // @[Mux.scala 31:69:@3507.4]
  wire [15:0] _T_6674; // @[Mux.scala 31:69:@3508.4]
  wire [15:0] _T_6675; // @[Mux.scala 31:69:@3509.4]
  wire [15:0] _T_6676; // @[Mux.scala 31:69:@3510.4]
  wire [15:0] _T_6677; // @[Mux.scala 31:69:@3511.4]
  wire [15:0] _T_6678; // @[Mux.scala 31:69:@3512.4]
  wire [15:0] _T_6679; // @[Mux.scala 31:69:@3513.4]
  wire [15:0] _T_6680; // @[Mux.scala 31:69:@3514.4]
  wire [15:0] _T_6681; // @[Mux.scala 31:69:@3515.4]
  wire [15:0] _T_6682; // @[Mux.scala 31:69:@3516.4]
  wire  _T_6683; // @[OneHot.scala 66:30:@3517.4]
  wire  _T_6684; // @[OneHot.scala 66:30:@3518.4]
  wire  _T_6685; // @[OneHot.scala 66:30:@3519.4]
  wire  _T_6686; // @[OneHot.scala 66:30:@3520.4]
  wire  _T_6687; // @[OneHot.scala 66:30:@3521.4]
  wire  _T_6688; // @[OneHot.scala 66:30:@3522.4]
  wire  _T_6689; // @[OneHot.scala 66:30:@3523.4]
  wire  _T_6690; // @[OneHot.scala 66:30:@3524.4]
  wire  _T_6691; // @[OneHot.scala 66:30:@3525.4]
  wire  _T_6692; // @[OneHot.scala 66:30:@3526.4]
  wire  _T_6693; // @[OneHot.scala 66:30:@3527.4]
  wire  _T_6694; // @[OneHot.scala 66:30:@3528.4]
  wire  _T_6695; // @[OneHot.scala 66:30:@3529.4]
  wire  _T_6696; // @[OneHot.scala 66:30:@3530.4]
  wire  _T_6697; // @[OneHot.scala 66:30:@3531.4]
  wire  _T_6698; // @[OneHot.scala 66:30:@3532.4]
  wire [15:0] _T_6739; // @[Mux.scala 31:69:@3550.4]
  wire [15:0] _T_6740; // @[Mux.scala 31:69:@3551.4]
  wire [15:0] _T_6741; // @[Mux.scala 31:69:@3552.4]
  wire [15:0] _T_6742; // @[Mux.scala 31:69:@3553.4]
  wire [15:0] _T_6743; // @[Mux.scala 31:69:@3554.4]
  wire [15:0] _T_6744; // @[Mux.scala 31:69:@3555.4]
  wire [15:0] _T_6745; // @[Mux.scala 31:69:@3556.4]
  wire [15:0] _T_6746; // @[Mux.scala 31:69:@3557.4]
  wire [15:0] _T_6747; // @[Mux.scala 31:69:@3558.4]
  wire [15:0] _T_6748; // @[Mux.scala 31:69:@3559.4]
  wire [15:0] _T_6749; // @[Mux.scala 31:69:@3560.4]
  wire [15:0] _T_6750; // @[Mux.scala 31:69:@3561.4]
  wire [15:0] _T_6751; // @[Mux.scala 31:69:@3562.4]
  wire [15:0] _T_6752; // @[Mux.scala 31:69:@3563.4]
  wire [15:0] _T_6753; // @[Mux.scala 31:69:@3564.4]
  wire [15:0] _T_6754; // @[Mux.scala 31:69:@3565.4]
  wire  _T_6755; // @[OneHot.scala 66:30:@3566.4]
  wire  _T_6756; // @[OneHot.scala 66:30:@3567.4]
  wire  _T_6757; // @[OneHot.scala 66:30:@3568.4]
  wire  _T_6758; // @[OneHot.scala 66:30:@3569.4]
  wire  _T_6759; // @[OneHot.scala 66:30:@3570.4]
  wire  _T_6760; // @[OneHot.scala 66:30:@3571.4]
  wire  _T_6761; // @[OneHot.scala 66:30:@3572.4]
  wire  _T_6762; // @[OneHot.scala 66:30:@3573.4]
  wire  _T_6763; // @[OneHot.scala 66:30:@3574.4]
  wire  _T_6764; // @[OneHot.scala 66:30:@3575.4]
  wire  _T_6765; // @[OneHot.scala 66:30:@3576.4]
  wire  _T_6766; // @[OneHot.scala 66:30:@3577.4]
  wire  _T_6767; // @[OneHot.scala 66:30:@3578.4]
  wire  _T_6768; // @[OneHot.scala 66:30:@3579.4]
  wire  _T_6769; // @[OneHot.scala 66:30:@3580.4]
  wire  _T_6770; // @[OneHot.scala 66:30:@3581.4]
  wire [15:0] _T_6811; // @[Mux.scala 31:69:@3599.4]
  wire [15:0] _T_6812; // @[Mux.scala 31:69:@3600.4]
  wire [15:0] _T_6813; // @[Mux.scala 31:69:@3601.4]
  wire [15:0] _T_6814; // @[Mux.scala 31:69:@3602.4]
  wire [15:0] _T_6815; // @[Mux.scala 31:69:@3603.4]
  wire [15:0] _T_6816; // @[Mux.scala 31:69:@3604.4]
  wire [15:0] _T_6817; // @[Mux.scala 31:69:@3605.4]
  wire [15:0] _T_6818; // @[Mux.scala 31:69:@3606.4]
  wire [15:0] _T_6819; // @[Mux.scala 31:69:@3607.4]
  wire [15:0] _T_6820; // @[Mux.scala 31:69:@3608.4]
  wire [15:0] _T_6821; // @[Mux.scala 31:69:@3609.4]
  wire [15:0] _T_6822; // @[Mux.scala 31:69:@3610.4]
  wire [15:0] _T_6823; // @[Mux.scala 31:69:@3611.4]
  wire [15:0] _T_6824; // @[Mux.scala 31:69:@3612.4]
  wire [15:0] _T_6825; // @[Mux.scala 31:69:@3613.4]
  wire [15:0] _T_6826; // @[Mux.scala 31:69:@3614.4]
  wire  _T_6827; // @[OneHot.scala 66:30:@3615.4]
  wire  _T_6828; // @[OneHot.scala 66:30:@3616.4]
  wire  _T_6829; // @[OneHot.scala 66:30:@3617.4]
  wire  _T_6830; // @[OneHot.scala 66:30:@3618.4]
  wire  _T_6831; // @[OneHot.scala 66:30:@3619.4]
  wire  _T_6832; // @[OneHot.scala 66:30:@3620.4]
  wire  _T_6833; // @[OneHot.scala 66:30:@3621.4]
  wire  _T_6834; // @[OneHot.scala 66:30:@3622.4]
  wire  _T_6835; // @[OneHot.scala 66:30:@3623.4]
  wire  _T_6836; // @[OneHot.scala 66:30:@3624.4]
  wire  _T_6837; // @[OneHot.scala 66:30:@3625.4]
  wire  _T_6838; // @[OneHot.scala 66:30:@3626.4]
  wire  _T_6839; // @[OneHot.scala 66:30:@3627.4]
  wire  _T_6840; // @[OneHot.scala 66:30:@3628.4]
  wire  _T_6841; // @[OneHot.scala 66:30:@3629.4]
  wire  _T_6842; // @[OneHot.scala 66:30:@3630.4]
  wire [15:0] _T_6883; // @[Mux.scala 31:69:@3648.4]
  wire [15:0] _T_6884; // @[Mux.scala 31:69:@3649.4]
  wire [15:0] _T_6885; // @[Mux.scala 31:69:@3650.4]
  wire [15:0] _T_6886; // @[Mux.scala 31:69:@3651.4]
  wire [15:0] _T_6887; // @[Mux.scala 31:69:@3652.4]
  wire [15:0] _T_6888; // @[Mux.scala 31:69:@3653.4]
  wire [15:0] _T_6889; // @[Mux.scala 31:69:@3654.4]
  wire [15:0] _T_6890; // @[Mux.scala 31:69:@3655.4]
  wire [15:0] _T_6891; // @[Mux.scala 31:69:@3656.4]
  wire [15:0] _T_6892; // @[Mux.scala 31:69:@3657.4]
  wire [15:0] _T_6893; // @[Mux.scala 31:69:@3658.4]
  wire [15:0] _T_6894; // @[Mux.scala 31:69:@3659.4]
  wire [15:0] _T_6895; // @[Mux.scala 31:69:@3660.4]
  wire [15:0] _T_6896; // @[Mux.scala 31:69:@3661.4]
  wire [15:0] _T_6897; // @[Mux.scala 31:69:@3662.4]
  wire [15:0] _T_6898; // @[Mux.scala 31:69:@3663.4]
  wire  _T_6899; // @[OneHot.scala 66:30:@3664.4]
  wire  _T_6900; // @[OneHot.scala 66:30:@3665.4]
  wire  _T_6901; // @[OneHot.scala 66:30:@3666.4]
  wire  _T_6902; // @[OneHot.scala 66:30:@3667.4]
  wire  _T_6903; // @[OneHot.scala 66:30:@3668.4]
  wire  _T_6904; // @[OneHot.scala 66:30:@3669.4]
  wire  _T_6905; // @[OneHot.scala 66:30:@3670.4]
  wire  _T_6906; // @[OneHot.scala 66:30:@3671.4]
  wire  _T_6907; // @[OneHot.scala 66:30:@3672.4]
  wire  _T_6908; // @[OneHot.scala 66:30:@3673.4]
  wire  _T_6909; // @[OneHot.scala 66:30:@3674.4]
  wire  _T_6910; // @[OneHot.scala 66:30:@3675.4]
  wire  _T_6911; // @[OneHot.scala 66:30:@3676.4]
  wire  _T_6912; // @[OneHot.scala 66:30:@3677.4]
  wire  _T_6913; // @[OneHot.scala 66:30:@3678.4]
  wire  _T_6914; // @[OneHot.scala 66:30:@3679.4]
  wire [15:0] _T_6955; // @[Mux.scala 31:69:@3697.4]
  wire [15:0] _T_6956; // @[Mux.scala 31:69:@3698.4]
  wire [15:0] _T_6957; // @[Mux.scala 31:69:@3699.4]
  wire [15:0] _T_6958; // @[Mux.scala 31:69:@3700.4]
  wire [15:0] _T_6959; // @[Mux.scala 31:69:@3701.4]
  wire [15:0] _T_6960; // @[Mux.scala 31:69:@3702.4]
  wire [15:0] _T_6961; // @[Mux.scala 31:69:@3703.4]
  wire [15:0] _T_6962; // @[Mux.scala 31:69:@3704.4]
  wire [15:0] _T_6963; // @[Mux.scala 31:69:@3705.4]
  wire [15:0] _T_6964; // @[Mux.scala 31:69:@3706.4]
  wire [15:0] _T_6965; // @[Mux.scala 31:69:@3707.4]
  wire [15:0] _T_6966; // @[Mux.scala 31:69:@3708.4]
  wire [15:0] _T_6967; // @[Mux.scala 31:69:@3709.4]
  wire [15:0] _T_6968; // @[Mux.scala 31:69:@3710.4]
  wire [15:0] _T_6969; // @[Mux.scala 31:69:@3711.4]
  wire [15:0] _T_6970; // @[Mux.scala 31:69:@3712.4]
  wire  _T_6971; // @[OneHot.scala 66:30:@3713.4]
  wire  _T_6972; // @[OneHot.scala 66:30:@3714.4]
  wire  _T_6973; // @[OneHot.scala 66:30:@3715.4]
  wire  _T_6974; // @[OneHot.scala 66:30:@3716.4]
  wire  _T_6975; // @[OneHot.scala 66:30:@3717.4]
  wire  _T_6976; // @[OneHot.scala 66:30:@3718.4]
  wire  _T_6977; // @[OneHot.scala 66:30:@3719.4]
  wire  _T_6978; // @[OneHot.scala 66:30:@3720.4]
  wire  _T_6979; // @[OneHot.scala 66:30:@3721.4]
  wire  _T_6980; // @[OneHot.scala 66:30:@3722.4]
  wire  _T_6981; // @[OneHot.scala 66:30:@3723.4]
  wire  _T_6982; // @[OneHot.scala 66:30:@3724.4]
  wire  _T_6983; // @[OneHot.scala 66:30:@3725.4]
  wire  _T_6984; // @[OneHot.scala 66:30:@3726.4]
  wire  _T_6985; // @[OneHot.scala 66:30:@3727.4]
  wire  _T_6986; // @[OneHot.scala 66:30:@3728.4]
  wire [15:0] _T_7027; // @[Mux.scala 31:69:@3746.4]
  wire [15:0] _T_7028; // @[Mux.scala 31:69:@3747.4]
  wire [15:0] _T_7029; // @[Mux.scala 31:69:@3748.4]
  wire [15:0] _T_7030; // @[Mux.scala 31:69:@3749.4]
  wire [15:0] _T_7031; // @[Mux.scala 31:69:@3750.4]
  wire [15:0] _T_7032; // @[Mux.scala 31:69:@3751.4]
  wire [15:0] _T_7033; // @[Mux.scala 31:69:@3752.4]
  wire [15:0] _T_7034; // @[Mux.scala 31:69:@3753.4]
  wire [15:0] _T_7035; // @[Mux.scala 31:69:@3754.4]
  wire [15:0] _T_7036; // @[Mux.scala 31:69:@3755.4]
  wire [15:0] _T_7037; // @[Mux.scala 31:69:@3756.4]
  wire [15:0] _T_7038; // @[Mux.scala 31:69:@3757.4]
  wire [15:0] _T_7039; // @[Mux.scala 31:69:@3758.4]
  wire [15:0] _T_7040; // @[Mux.scala 31:69:@3759.4]
  wire [15:0] _T_7041; // @[Mux.scala 31:69:@3760.4]
  wire [15:0] _T_7042; // @[Mux.scala 31:69:@3761.4]
  wire  _T_7043; // @[OneHot.scala 66:30:@3762.4]
  wire  _T_7044; // @[OneHot.scala 66:30:@3763.4]
  wire  _T_7045; // @[OneHot.scala 66:30:@3764.4]
  wire  _T_7046; // @[OneHot.scala 66:30:@3765.4]
  wire  _T_7047; // @[OneHot.scala 66:30:@3766.4]
  wire  _T_7048; // @[OneHot.scala 66:30:@3767.4]
  wire  _T_7049; // @[OneHot.scala 66:30:@3768.4]
  wire  _T_7050; // @[OneHot.scala 66:30:@3769.4]
  wire  _T_7051; // @[OneHot.scala 66:30:@3770.4]
  wire  _T_7052; // @[OneHot.scala 66:30:@3771.4]
  wire  _T_7053; // @[OneHot.scala 66:30:@3772.4]
  wire  _T_7054; // @[OneHot.scala 66:30:@3773.4]
  wire  _T_7055; // @[OneHot.scala 66:30:@3774.4]
  wire  _T_7056; // @[OneHot.scala 66:30:@3775.4]
  wire  _T_7057; // @[OneHot.scala 66:30:@3776.4]
  wire  _T_7058; // @[OneHot.scala 66:30:@3777.4]
  wire [15:0] _T_7099; // @[Mux.scala 31:69:@3795.4]
  wire [15:0] _T_7100; // @[Mux.scala 31:69:@3796.4]
  wire [15:0] _T_7101; // @[Mux.scala 31:69:@3797.4]
  wire [15:0] _T_7102; // @[Mux.scala 31:69:@3798.4]
  wire [15:0] _T_7103; // @[Mux.scala 31:69:@3799.4]
  wire [15:0] _T_7104; // @[Mux.scala 31:69:@3800.4]
  wire [15:0] _T_7105; // @[Mux.scala 31:69:@3801.4]
  wire [15:0] _T_7106; // @[Mux.scala 31:69:@3802.4]
  wire [15:0] _T_7107; // @[Mux.scala 31:69:@3803.4]
  wire [15:0] _T_7108; // @[Mux.scala 31:69:@3804.4]
  wire [15:0] _T_7109; // @[Mux.scala 31:69:@3805.4]
  wire [15:0] _T_7110; // @[Mux.scala 31:69:@3806.4]
  wire [15:0] _T_7111; // @[Mux.scala 31:69:@3807.4]
  wire [15:0] _T_7112; // @[Mux.scala 31:69:@3808.4]
  wire [15:0] _T_7113; // @[Mux.scala 31:69:@3809.4]
  wire [15:0] _T_7114; // @[Mux.scala 31:69:@3810.4]
  wire  _T_7115; // @[OneHot.scala 66:30:@3811.4]
  wire  _T_7116; // @[OneHot.scala 66:30:@3812.4]
  wire  _T_7117; // @[OneHot.scala 66:30:@3813.4]
  wire  _T_7118; // @[OneHot.scala 66:30:@3814.4]
  wire  _T_7119; // @[OneHot.scala 66:30:@3815.4]
  wire  _T_7120; // @[OneHot.scala 66:30:@3816.4]
  wire  _T_7121; // @[OneHot.scala 66:30:@3817.4]
  wire  _T_7122; // @[OneHot.scala 66:30:@3818.4]
  wire  _T_7123; // @[OneHot.scala 66:30:@3819.4]
  wire  _T_7124; // @[OneHot.scala 66:30:@3820.4]
  wire  _T_7125; // @[OneHot.scala 66:30:@3821.4]
  wire  _T_7126; // @[OneHot.scala 66:30:@3822.4]
  wire  _T_7127; // @[OneHot.scala 66:30:@3823.4]
  wire  _T_7128; // @[OneHot.scala 66:30:@3824.4]
  wire  _T_7129; // @[OneHot.scala 66:30:@3825.4]
  wire  _T_7130; // @[OneHot.scala 66:30:@3826.4]
  wire [15:0] _T_7171; // @[Mux.scala 31:69:@3844.4]
  wire [15:0] _T_7172; // @[Mux.scala 31:69:@3845.4]
  wire [15:0] _T_7173; // @[Mux.scala 31:69:@3846.4]
  wire [15:0] _T_7174; // @[Mux.scala 31:69:@3847.4]
  wire [15:0] _T_7175; // @[Mux.scala 31:69:@3848.4]
  wire [15:0] _T_7176; // @[Mux.scala 31:69:@3849.4]
  wire [15:0] _T_7177; // @[Mux.scala 31:69:@3850.4]
  wire [15:0] _T_7178; // @[Mux.scala 31:69:@3851.4]
  wire [15:0] _T_7179; // @[Mux.scala 31:69:@3852.4]
  wire [15:0] _T_7180; // @[Mux.scala 31:69:@3853.4]
  wire [15:0] _T_7181; // @[Mux.scala 31:69:@3854.4]
  wire [15:0] _T_7182; // @[Mux.scala 31:69:@3855.4]
  wire [15:0] _T_7183; // @[Mux.scala 31:69:@3856.4]
  wire [15:0] _T_7184; // @[Mux.scala 31:69:@3857.4]
  wire [15:0] _T_7185; // @[Mux.scala 31:69:@3858.4]
  wire [15:0] _T_7186; // @[Mux.scala 31:69:@3859.4]
  wire  _T_7187; // @[OneHot.scala 66:30:@3860.4]
  wire  _T_7188; // @[OneHot.scala 66:30:@3861.4]
  wire  _T_7189; // @[OneHot.scala 66:30:@3862.4]
  wire  _T_7190; // @[OneHot.scala 66:30:@3863.4]
  wire  _T_7191; // @[OneHot.scala 66:30:@3864.4]
  wire  _T_7192; // @[OneHot.scala 66:30:@3865.4]
  wire  _T_7193; // @[OneHot.scala 66:30:@3866.4]
  wire  _T_7194; // @[OneHot.scala 66:30:@3867.4]
  wire  _T_7195; // @[OneHot.scala 66:30:@3868.4]
  wire  _T_7196; // @[OneHot.scala 66:30:@3869.4]
  wire  _T_7197; // @[OneHot.scala 66:30:@3870.4]
  wire  _T_7198; // @[OneHot.scala 66:30:@3871.4]
  wire  _T_7199; // @[OneHot.scala 66:30:@3872.4]
  wire  _T_7200; // @[OneHot.scala 66:30:@3873.4]
  wire  _T_7201; // @[OneHot.scala 66:30:@3874.4]
  wire  _T_7202; // @[OneHot.scala 66:30:@3875.4]
  wire [15:0] _T_7243; // @[Mux.scala 31:69:@3893.4]
  wire [15:0] _T_7244; // @[Mux.scala 31:69:@3894.4]
  wire [15:0] _T_7245; // @[Mux.scala 31:69:@3895.4]
  wire [15:0] _T_7246; // @[Mux.scala 31:69:@3896.4]
  wire [15:0] _T_7247; // @[Mux.scala 31:69:@3897.4]
  wire [15:0] _T_7248; // @[Mux.scala 31:69:@3898.4]
  wire [15:0] _T_7249; // @[Mux.scala 31:69:@3899.4]
  wire [15:0] _T_7250; // @[Mux.scala 31:69:@3900.4]
  wire [15:0] _T_7251; // @[Mux.scala 31:69:@3901.4]
  wire [15:0] _T_7252; // @[Mux.scala 31:69:@3902.4]
  wire [15:0] _T_7253; // @[Mux.scala 31:69:@3903.4]
  wire [15:0] _T_7254; // @[Mux.scala 31:69:@3904.4]
  wire [15:0] _T_7255; // @[Mux.scala 31:69:@3905.4]
  wire [15:0] _T_7256; // @[Mux.scala 31:69:@3906.4]
  wire [15:0] _T_7257; // @[Mux.scala 31:69:@3907.4]
  wire [15:0] _T_7258; // @[Mux.scala 31:69:@3908.4]
  wire  _T_7259; // @[OneHot.scala 66:30:@3909.4]
  wire  _T_7260; // @[OneHot.scala 66:30:@3910.4]
  wire  _T_7261; // @[OneHot.scala 66:30:@3911.4]
  wire  _T_7262; // @[OneHot.scala 66:30:@3912.4]
  wire  _T_7263; // @[OneHot.scala 66:30:@3913.4]
  wire  _T_7264; // @[OneHot.scala 66:30:@3914.4]
  wire  _T_7265; // @[OneHot.scala 66:30:@3915.4]
  wire  _T_7266; // @[OneHot.scala 66:30:@3916.4]
  wire  _T_7267; // @[OneHot.scala 66:30:@3917.4]
  wire  _T_7268; // @[OneHot.scala 66:30:@3918.4]
  wire  _T_7269; // @[OneHot.scala 66:30:@3919.4]
  wire  _T_7270; // @[OneHot.scala 66:30:@3920.4]
  wire  _T_7271; // @[OneHot.scala 66:30:@3921.4]
  wire  _T_7272; // @[OneHot.scala 66:30:@3922.4]
  wire  _T_7273; // @[OneHot.scala 66:30:@3923.4]
  wire  _T_7274; // @[OneHot.scala 66:30:@3924.4]
  wire [15:0] _T_7315; // @[Mux.scala 31:69:@3942.4]
  wire [15:0] _T_7316; // @[Mux.scala 31:69:@3943.4]
  wire [15:0] _T_7317; // @[Mux.scala 31:69:@3944.4]
  wire [15:0] _T_7318; // @[Mux.scala 31:69:@3945.4]
  wire [15:0] _T_7319; // @[Mux.scala 31:69:@3946.4]
  wire [15:0] _T_7320; // @[Mux.scala 31:69:@3947.4]
  wire [15:0] _T_7321; // @[Mux.scala 31:69:@3948.4]
  wire [15:0] _T_7322; // @[Mux.scala 31:69:@3949.4]
  wire [15:0] _T_7323; // @[Mux.scala 31:69:@3950.4]
  wire [15:0] _T_7324; // @[Mux.scala 31:69:@3951.4]
  wire [15:0] _T_7325; // @[Mux.scala 31:69:@3952.4]
  wire [15:0] _T_7326; // @[Mux.scala 31:69:@3953.4]
  wire [15:0] _T_7327; // @[Mux.scala 31:69:@3954.4]
  wire [15:0] _T_7328; // @[Mux.scala 31:69:@3955.4]
  wire [15:0] _T_7329; // @[Mux.scala 31:69:@3956.4]
  wire [15:0] _T_7330; // @[Mux.scala 31:69:@3957.4]
  wire  _T_7331; // @[OneHot.scala 66:30:@3958.4]
  wire  _T_7332; // @[OneHot.scala 66:30:@3959.4]
  wire  _T_7333; // @[OneHot.scala 66:30:@3960.4]
  wire  _T_7334; // @[OneHot.scala 66:30:@3961.4]
  wire  _T_7335; // @[OneHot.scala 66:30:@3962.4]
  wire  _T_7336; // @[OneHot.scala 66:30:@3963.4]
  wire  _T_7337; // @[OneHot.scala 66:30:@3964.4]
  wire  _T_7338; // @[OneHot.scala 66:30:@3965.4]
  wire  _T_7339; // @[OneHot.scala 66:30:@3966.4]
  wire  _T_7340; // @[OneHot.scala 66:30:@3967.4]
  wire  _T_7341; // @[OneHot.scala 66:30:@3968.4]
  wire  _T_7342; // @[OneHot.scala 66:30:@3969.4]
  wire  _T_7343; // @[OneHot.scala 66:30:@3970.4]
  wire  _T_7344; // @[OneHot.scala 66:30:@3971.4]
  wire  _T_7345; // @[OneHot.scala 66:30:@3972.4]
  wire  _T_7346; // @[OneHot.scala 66:30:@3973.4]
  wire [7:0] _T_7411; // @[Mux.scala 19:72:@3997.4]
  wire [15:0] _T_7419; // @[Mux.scala 19:72:@4005.4]
  wire [15:0] _T_7421; // @[Mux.scala 19:72:@4006.4]
  wire [7:0] _T_7428; // @[Mux.scala 19:72:@4013.4]
  wire [15:0] _T_7436; // @[Mux.scala 19:72:@4021.4]
  wire [15:0] _T_7438; // @[Mux.scala 19:72:@4022.4]
  wire [7:0] _T_7445; // @[Mux.scala 19:72:@4029.4]
  wire [15:0] _T_7453; // @[Mux.scala 19:72:@4037.4]
  wire [15:0] _T_7455; // @[Mux.scala 19:72:@4038.4]
  wire [7:0] _T_7462; // @[Mux.scala 19:72:@4045.4]
  wire [15:0] _T_7470; // @[Mux.scala 19:72:@4053.4]
  wire [15:0] _T_7472; // @[Mux.scala 19:72:@4054.4]
  wire [7:0] _T_7479; // @[Mux.scala 19:72:@4061.4]
  wire [15:0] _T_7487; // @[Mux.scala 19:72:@4069.4]
  wire [15:0] _T_7489; // @[Mux.scala 19:72:@4070.4]
  wire [7:0] _T_7496; // @[Mux.scala 19:72:@4077.4]
  wire [15:0] _T_7504; // @[Mux.scala 19:72:@4085.4]
  wire [15:0] _T_7506; // @[Mux.scala 19:72:@4086.4]
  wire [7:0] _T_7513; // @[Mux.scala 19:72:@4093.4]
  wire [15:0] _T_7521; // @[Mux.scala 19:72:@4101.4]
  wire [15:0] _T_7523; // @[Mux.scala 19:72:@4102.4]
  wire [7:0] _T_7530; // @[Mux.scala 19:72:@4109.4]
  wire [15:0] _T_7538; // @[Mux.scala 19:72:@4117.4]
  wire [15:0] _T_7540; // @[Mux.scala 19:72:@4118.4]
  wire [7:0] _T_7547; // @[Mux.scala 19:72:@4125.4]
  wire [15:0] _T_7555; // @[Mux.scala 19:72:@4133.4]
  wire [15:0] _T_7557; // @[Mux.scala 19:72:@4134.4]
  wire [7:0] _T_7564; // @[Mux.scala 19:72:@4141.4]
  wire [15:0] _T_7572; // @[Mux.scala 19:72:@4149.4]
  wire [15:0] _T_7574; // @[Mux.scala 19:72:@4150.4]
  wire [7:0] _T_7581; // @[Mux.scala 19:72:@4157.4]
  wire [15:0] _T_7589; // @[Mux.scala 19:72:@4165.4]
  wire [15:0] _T_7591; // @[Mux.scala 19:72:@4166.4]
  wire [7:0] _T_7598; // @[Mux.scala 19:72:@4173.4]
  wire [15:0] _T_7606; // @[Mux.scala 19:72:@4181.4]
  wire [15:0] _T_7608; // @[Mux.scala 19:72:@4182.4]
  wire [7:0] _T_7615; // @[Mux.scala 19:72:@4189.4]
  wire [15:0] _T_7623; // @[Mux.scala 19:72:@4197.4]
  wire [15:0] _T_7625; // @[Mux.scala 19:72:@4198.4]
  wire [7:0] _T_7632; // @[Mux.scala 19:72:@4205.4]
  wire [15:0] _T_7640; // @[Mux.scala 19:72:@4213.4]
  wire [15:0] _T_7642; // @[Mux.scala 19:72:@4214.4]
  wire [7:0] _T_7649; // @[Mux.scala 19:72:@4221.4]
  wire [15:0] _T_7657; // @[Mux.scala 19:72:@4229.4]
  wire [15:0] _T_7659; // @[Mux.scala 19:72:@4230.4]
  wire [7:0] _T_7666; // @[Mux.scala 19:72:@4237.4]
  wire [15:0] _T_7674; // @[Mux.scala 19:72:@4245.4]
  wire [15:0] _T_7676; // @[Mux.scala 19:72:@4246.4]
  wire [15:0] _T_7677; // @[Mux.scala 19:72:@4247.4]
  wire [15:0] _T_7678; // @[Mux.scala 19:72:@4248.4]
  wire [15:0] _T_7679; // @[Mux.scala 19:72:@4249.4]
  wire [15:0] _T_7680; // @[Mux.scala 19:72:@4250.4]
  wire [15:0] _T_7681; // @[Mux.scala 19:72:@4251.4]
  wire [15:0] _T_7682; // @[Mux.scala 19:72:@4252.4]
  wire [15:0] _T_7683; // @[Mux.scala 19:72:@4253.4]
  wire [15:0] _T_7684; // @[Mux.scala 19:72:@4254.4]
  wire [15:0] _T_7685; // @[Mux.scala 19:72:@4255.4]
  wire [15:0] _T_7686; // @[Mux.scala 19:72:@4256.4]
  wire [15:0] _T_7687; // @[Mux.scala 19:72:@4257.4]
  wire [15:0] _T_7688; // @[Mux.scala 19:72:@4258.4]
  wire [15:0] _T_7689; // @[Mux.scala 19:72:@4259.4]
  wire [15:0] _T_7690; // @[Mux.scala 19:72:@4260.4]
  wire [15:0] _T_7691; // @[Mux.scala 19:72:@4261.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@4265.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@4267.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@4269.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@4271.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@4273.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@4275.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@4277.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@4279.4]
  wire  inputDataPriorityPorts_0_8; // @[Mux.scala 19:72:@4281.4]
  wire  inputDataPriorityPorts_0_9; // @[Mux.scala 19:72:@4283.4]
  wire  inputDataPriorityPorts_0_10; // @[Mux.scala 19:72:@4285.4]
  wire  inputDataPriorityPorts_0_11; // @[Mux.scala 19:72:@4287.4]
  wire  inputDataPriorityPorts_0_12; // @[Mux.scala 19:72:@4289.4]
  wire  inputDataPriorityPorts_0_13; // @[Mux.scala 19:72:@4291.4]
  wire  inputDataPriorityPorts_0_14; // @[Mux.scala 19:72:@4293.4]
  wire  inputDataPriorityPorts_0_15; // @[Mux.scala 19:72:@4295.4]
  wire  _T_7835; // @[StoreQueue.scala 192:88:@4314.4]
  wire  _T_7838; // @[StoreQueue.scala 192:88:@4316.4]
  wire  _T_7841; // @[StoreQueue.scala 192:88:@4318.4]
  wire  _T_7844; // @[StoreQueue.scala 192:88:@4320.4]
  wire  _T_7847; // @[StoreQueue.scala 192:88:@4322.4]
  wire  _T_7850; // @[StoreQueue.scala 192:88:@4324.4]
  wire  _T_7853; // @[StoreQueue.scala 192:88:@4326.4]
  wire  _T_7856; // @[StoreQueue.scala 192:88:@4328.4]
  wire  _T_7859; // @[StoreQueue.scala 192:88:@4330.4]
  wire  _T_7862; // @[StoreQueue.scala 192:88:@4332.4]
  wire  _T_7865; // @[StoreQueue.scala 192:88:@4334.4]
  wire  _T_7868; // @[StoreQueue.scala 192:88:@4336.4]
  wire  _T_7871; // @[StoreQueue.scala 192:88:@4338.4]
  wire  _T_7874; // @[StoreQueue.scala 192:88:@4340.4]
  wire  _T_7877; // @[StoreQueue.scala 192:88:@4342.4]
  wire  _T_7880; // @[StoreQueue.scala 192:88:@4344.4]
  wire  _T_7905; // @[StoreQueue.scala 193:88:@4363.4]
  wire  _T_7908; // @[StoreQueue.scala 193:88:@4365.4]
  wire  _T_7911; // @[StoreQueue.scala 193:88:@4367.4]
  wire  _T_7914; // @[StoreQueue.scala 193:88:@4369.4]
  wire  _T_7917; // @[StoreQueue.scala 193:88:@4371.4]
  wire  _T_7920; // @[StoreQueue.scala 193:88:@4373.4]
  wire  _T_7923; // @[StoreQueue.scala 193:88:@4375.4]
  wire  _T_7926; // @[StoreQueue.scala 193:88:@4377.4]
  wire  _T_7929; // @[StoreQueue.scala 193:88:@4379.4]
  wire  _T_7932; // @[StoreQueue.scala 193:88:@4381.4]
  wire  _T_7935; // @[StoreQueue.scala 193:88:@4383.4]
  wire  _T_7938; // @[StoreQueue.scala 193:88:@4385.4]
  wire  _T_7941; // @[StoreQueue.scala 193:88:@4387.4]
  wire  _T_7944; // @[StoreQueue.scala 193:88:@4389.4]
  wire  _T_7947; // @[StoreQueue.scala 193:88:@4391.4]
  wire  _T_7950; // @[StoreQueue.scala 193:88:@4393.4]
  wire [15:0] _T_8033; // @[Mux.scala 31:69:@4447.4]
  wire [15:0] _T_8034; // @[Mux.scala 31:69:@4448.4]
  wire [15:0] _T_8035; // @[Mux.scala 31:69:@4449.4]
  wire [15:0] _T_8036; // @[Mux.scala 31:69:@4450.4]
  wire [15:0] _T_8037; // @[Mux.scala 31:69:@4451.4]
  wire [15:0] _T_8038; // @[Mux.scala 31:69:@4452.4]
  wire [15:0] _T_8039; // @[Mux.scala 31:69:@4453.4]
  wire [15:0] _T_8040; // @[Mux.scala 31:69:@4454.4]
  wire [15:0] _T_8041; // @[Mux.scala 31:69:@4455.4]
  wire [15:0] _T_8042; // @[Mux.scala 31:69:@4456.4]
  wire [15:0] _T_8043; // @[Mux.scala 31:69:@4457.4]
  wire [15:0] _T_8044; // @[Mux.scala 31:69:@4458.4]
  wire [15:0] _T_8045; // @[Mux.scala 31:69:@4459.4]
  wire [15:0] _T_8046; // @[Mux.scala 31:69:@4460.4]
  wire [15:0] _T_8047; // @[Mux.scala 31:69:@4461.4]
  wire [15:0] _T_8048; // @[Mux.scala 31:69:@4462.4]
  wire  _T_8049; // @[OneHot.scala 66:30:@4463.4]
  wire  _T_8050; // @[OneHot.scala 66:30:@4464.4]
  wire  _T_8051; // @[OneHot.scala 66:30:@4465.4]
  wire  _T_8052; // @[OneHot.scala 66:30:@4466.4]
  wire  _T_8053; // @[OneHot.scala 66:30:@4467.4]
  wire  _T_8054; // @[OneHot.scala 66:30:@4468.4]
  wire  _T_8055; // @[OneHot.scala 66:30:@4469.4]
  wire  _T_8056; // @[OneHot.scala 66:30:@4470.4]
  wire  _T_8057; // @[OneHot.scala 66:30:@4471.4]
  wire  _T_8058; // @[OneHot.scala 66:30:@4472.4]
  wire  _T_8059; // @[OneHot.scala 66:30:@4473.4]
  wire  _T_8060; // @[OneHot.scala 66:30:@4474.4]
  wire  _T_8061; // @[OneHot.scala 66:30:@4475.4]
  wire  _T_8062; // @[OneHot.scala 66:30:@4476.4]
  wire  _T_8063; // @[OneHot.scala 66:30:@4477.4]
  wire  _T_8064; // @[OneHot.scala 66:30:@4478.4]
  wire [15:0] _T_8105; // @[Mux.scala 31:69:@4496.4]
  wire [15:0] _T_8106; // @[Mux.scala 31:69:@4497.4]
  wire [15:0] _T_8107; // @[Mux.scala 31:69:@4498.4]
  wire [15:0] _T_8108; // @[Mux.scala 31:69:@4499.4]
  wire [15:0] _T_8109; // @[Mux.scala 31:69:@4500.4]
  wire [15:0] _T_8110; // @[Mux.scala 31:69:@4501.4]
  wire [15:0] _T_8111; // @[Mux.scala 31:69:@4502.4]
  wire [15:0] _T_8112; // @[Mux.scala 31:69:@4503.4]
  wire [15:0] _T_8113; // @[Mux.scala 31:69:@4504.4]
  wire [15:0] _T_8114; // @[Mux.scala 31:69:@4505.4]
  wire [15:0] _T_8115; // @[Mux.scala 31:69:@4506.4]
  wire [15:0] _T_8116; // @[Mux.scala 31:69:@4507.4]
  wire [15:0] _T_8117; // @[Mux.scala 31:69:@4508.4]
  wire [15:0] _T_8118; // @[Mux.scala 31:69:@4509.4]
  wire [15:0] _T_8119; // @[Mux.scala 31:69:@4510.4]
  wire [15:0] _T_8120; // @[Mux.scala 31:69:@4511.4]
  wire  _T_8121; // @[OneHot.scala 66:30:@4512.4]
  wire  _T_8122; // @[OneHot.scala 66:30:@4513.4]
  wire  _T_8123; // @[OneHot.scala 66:30:@4514.4]
  wire  _T_8124; // @[OneHot.scala 66:30:@4515.4]
  wire  _T_8125; // @[OneHot.scala 66:30:@4516.4]
  wire  _T_8126; // @[OneHot.scala 66:30:@4517.4]
  wire  _T_8127; // @[OneHot.scala 66:30:@4518.4]
  wire  _T_8128; // @[OneHot.scala 66:30:@4519.4]
  wire  _T_8129; // @[OneHot.scala 66:30:@4520.4]
  wire  _T_8130; // @[OneHot.scala 66:30:@4521.4]
  wire  _T_8131; // @[OneHot.scala 66:30:@4522.4]
  wire  _T_8132; // @[OneHot.scala 66:30:@4523.4]
  wire  _T_8133; // @[OneHot.scala 66:30:@4524.4]
  wire  _T_8134; // @[OneHot.scala 66:30:@4525.4]
  wire  _T_8135; // @[OneHot.scala 66:30:@4526.4]
  wire  _T_8136; // @[OneHot.scala 66:30:@4527.4]
  wire [15:0] _T_8177; // @[Mux.scala 31:69:@4545.4]
  wire [15:0] _T_8178; // @[Mux.scala 31:69:@4546.4]
  wire [15:0] _T_8179; // @[Mux.scala 31:69:@4547.4]
  wire [15:0] _T_8180; // @[Mux.scala 31:69:@4548.4]
  wire [15:0] _T_8181; // @[Mux.scala 31:69:@4549.4]
  wire [15:0] _T_8182; // @[Mux.scala 31:69:@4550.4]
  wire [15:0] _T_8183; // @[Mux.scala 31:69:@4551.4]
  wire [15:0] _T_8184; // @[Mux.scala 31:69:@4552.4]
  wire [15:0] _T_8185; // @[Mux.scala 31:69:@4553.4]
  wire [15:0] _T_8186; // @[Mux.scala 31:69:@4554.4]
  wire [15:0] _T_8187; // @[Mux.scala 31:69:@4555.4]
  wire [15:0] _T_8188; // @[Mux.scala 31:69:@4556.4]
  wire [15:0] _T_8189; // @[Mux.scala 31:69:@4557.4]
  wire [15:0] _T_8190; // @[Mux.scala 31:69:@4558.4]
  wire [15:0] _T_8191; // @[Mux.scala 31:69:@4559.4]
  wire [15:0] _T_8192; // @[Mux.scala 31:69:@4560.4]
  wire  _T_8193; // @[OneHot.scala 66:30:@4561.4]
  wire  _T_8194; // @[OneHot.scala 66:30:@4562.4]
  wire  _T_8195; // @[OneHot.scala 66:30:@4563.4]
  wire  _T_8196; // @[OneHot.scala 66:30:@4564.4]
  wire  _T_8197; // @[OneHot.scala 66:30:@4565.4]
  wire  _T_8198; // @[OneHot.scala 66:30:@4566.4]
  wire  _T_8199; // @[OneHot.scala 66:30:@4567.4]
  wire  _T_8200; // @[OneHot.scala 66:30:@4568.4]
  wire  _T_8201; // @[OneHot.scala 66:30:@4569.4]
  wire  _T_8202; // @[OneHot.scala 66:30:@4570.4]
  wire  _T_8203; // @[OneHot.scala 66:30:@4571.4]
  wire  _T_8204; // @[OneHot.scala 66:30:@4572.4]
  wire  _T_8205; // @[OneHot.scala 66:30:@4573.4]
  wire  _T_8206; // @[OneHot.scala 66:30:@4574.4]
  wire  _T_8207; // @[OneHot.scala 66:30:@4575.4]
  wire  _T_8208; // @[OneHot.scala 66:30:@4576.4]
  wire [15:0] _T_8249; // @[Mux.scala 31:69:@4594.4]
  wire [15:0] _T_8250; // @[Mux.scala 31:69:@4595.4]
  wire [15:0] _T_8251; // @[Mux.scala 31:69:@4596.4]
  wire [15:0] _T_8252; // @[Mux.scala 31:69:@4597.4]
  wire [15:0] _T_8253; // @[Mux.scala 31:69:@4598.4]
  wire [15:0] _T_8254; // @[Mux.scala 31:69:@4599.4]
  wire [15:0] _T_8255; // @[Mux.scala 31:69:@4600.4]
  wire [15:0] _T_8256; // @[Mux.scala 31:69:@4601.4]
  wire [15:0] _T_8257; // @[Mux.scala 31:69:@4602.4]
  wire [15:0] _T_8258; // @[Mux.scala 31:69:@4603.4]
  wire [15:0] _T_8259; // @[Mux.scala 31:69:@4604.4]
  wire [15:0] _T_8260; // @[Mux.scala 31:69:@4605.4]
  wire [15:0] _T_8261; // @[Mux.scala 31:69:@4606.4]
  wire [15:0] _T_8262; // @[Mux.scala 31:69:@4607.4]
  wire [15:0] _T_8263; // @[Mux.scala 31:69:@4608.4]
  wire [15:0] _T_8264; // @[Mux.scala 31:69:@4609.4]
  wire  _T_8265; // @[OneHot.scala 66:30:@4610.4]
  wire  _T_8266; // @[OneHot.scala 66:30:@4611.4]
  wire  _T_8267; // @[OneHot.scala 66:30:@4612.4]
  wire  _T_8268; // @[OneHot.scala 66:30:@4613.4]
  wire  _T_8269; // @[OneHot.scala 66:30:@4614.4]
  wire  _T_8270; // @[OneHot.scala 66:30:@4615.4]
  wire  _T_8271; // @[OneHot.scala 66:30:@4616.4]
  wire  _T_8272; // @[OneHot.scala 66:30:@4617.4]
  wire  _T_8273; // @[OneHot.scala 66:30:@4618.4]
  wire  _T_8274; // @[OneHot.scala 66:30:@4619.4]
  wire  _T_8275; // @[OneHot.scala 66:30:@4620.4]
  wire  _T_8276; // @[OneHot.scala 66:30:@4621.4]
  wire  _T_8277; // @[OneHot.scala 66:30:@4622.4]
  wire  _T_8278; // @[OneHot.scala 66:30:@4623.4]
  wire  _T_8279; // @[OneHot.scala 66:30:@4624.4]
  wire  _T_8280; // @[OneHot.scala 66:30:@4625.4]
  wire [15:0] _T_8321; // @[Mux.scala 31:69:@4643.4]
  wire [15:0] _T_8322; // @[Mux.scala 31:69:@4644.4]
  wire [15:0] _T_8323; // @[Mux.scala 31:69:@4645.4]
  wire [15:0] _T_8324; // @[Mux.scala 31:69:@4646.4]
  wire [15:0] _T_8325; // @[Mux.scala 31:69:@4647.4]
  wire [15:0] _T_8326; // @[Mux.scala 31:69:@4648.4]
  wire [15:0] _T_8327; // @[Mux.scala 31:69:@4649.4]
  wire [15:0] _T_8328; // @[Mux.scala 31:69:@4650.4]
  wire [15:0] _T_8329; // @[Mux.scala 31:69:@4651.4]
  wire [15:0] _T_8330; // @[Mux.scala 31:69:@4652.4]
  wire [15:0] _T_8331; // @[Mux.scala 31:69:@4653.4]
  wire [15:0] _T_8332; // @[Mux.scala 31:69:@4654.4]
  wire [15:0] _T_8333; // @[Mux.scala 31:69:@4655.4]
  wire [15:0] _T_8334; // @[Mux.scala 31:69:@4656.4]
  wire [15:0] _T_8335; // @[Mux.scala 31:69:@4657.4]
  wire [15:0] _T_8336; // @[Mux.scala 31:69:@4658.4]
  wire  _T_8337; // @[OneHot.scala 66:30:@4659.4]
  wire  _T_8338; // @[OneHot.scala 66:30:@4660.4]
  wire  _T_8339; // @[OneHot.scala 66:30:@4661.4]
  wire  _T_8340; // @[OneHot.scala 66:30:@4662.4]
  wire  _T_8341; // @[OneHot.scala 66:30:@4663.4]
  wire  _T_8342; // @[OneHot.scala 66:30:@4664.4]
  wire  _T_8343; // @[OneHot.scala 66:30:@4665.4]
  wire  _T_8344; // @[OneHot.scala 66:30:@4666.4]
  wire  _T_8345; // @[OneHot.scala 66:30:@4667.4]
  wire  _T_8346; // @[OneHot.scala 66:30:@4668.4]
  wire  _T_8347; // @[OneHot.scala 66:30:@4669.4]
  wire  _T_8348; // @[OneHot.scala 66:30:@4670.4]
  wire  _T_8349; // @[OneHot.scala 66:30:@4671.4]
  wire  _T_8350; // @[OneHot.scala 66:30:@4672.4]
  wire  _T_8351; // @[OneHot.scala 66:30:@4673.4]
  wire  _T_8352; // @[OneHot.scala 66:30:@4674.4]
  wire [15:0] _T_8393; // @[Mux.scala 31:69:@4692.4]
  wire [15:0] _T_8394; // @[Mux.scala 31:69:@4693.4]
  wire [15:0] _T_8395; // @[Mux.scala 31:69:@4694.4]
  wire [15:0] _T_8396; // @[Mux.scala 31:69:@4695.4]
  wire [15:0] _T_8397; // @[Mux.scala 31:69:@4696.4]
  wire [15:0] _T_8398; // @[Mux.scala 31:69:@4697.4]
  wire [15:0] _T_8399; // @[Mux.scala 31:69:@4698.4]
  wire [15:0] _T_8400; // @[Mux.scala 31:69:@4699.4]
  wire [15:0] _T_8401; // @[Mux.scala 31:69:@4700.4]
  wire [15:0] _T_8402; // @[Mux.scala 31:69:@4701.4]
  wire [15:0] _T_8403; // @[Mux.scala 31:69:@4702.4]
  wire [15:0] _T_8404; // @[Mux.scala 31:69:@4703.4]
  wire [15:0] _T_8405; // @[Mux.scala 31:69:@4704.4]
  wire [15:0] _T_8406; // @[Mux.scala 31:69:@4705.4]
  wire [15:0] _T_8407; // @[Mux.scala 31:69:@4706.4]
  wire [15:0] _T_8408; // @[Mux.scala 31:69:@4707.4]
  wire  _T_8409; // @[OneHot.scala 66:30:@4708.4]
  wire  _T_8410; // @[OneHot.scala 66:30:@4709.4]
  wire  _T_8411; // @[OneHot.scala 66:30:@4710.4]
  wire  _T_8412; // @[OneHot.scala 66:30:@4711.4]
  wire  _T_8413; // @[OneHot.scala 66:30:@4712.4]
  wire  _T_8414; // @[OneHot.scala 66:30:@4713.4]
  wire  _T_8415; // @[OneHot.scala 66:30:@4714.4]
  wire  _T_8416; // @[OneHot.scala 66:30:@4715.4]
  wire  _T_8417; // @[OneHot.scala 66:30:@4716.4]
  wire  _T_8418; // @[OneHot.scala 66:30:@4717.4]
  wire  _T_8419; // @[OneHot.scala 66:30:@4718.4]
  wire  _T_8420; // @[OneHot.scala 66:30:@4719.4]
  wire  _T_8421; // @[OneHot.scala 66:30:@4720.4]
  wire  _T_8422; // @[OneHot.scala 66:30:@4721.4]
  wire  _T_8423; // @[OneHot.scala 66:30:@4722.4]
  wire  _T_8424; // @[OneHot.scala 66:30:@4723.4]
  wire [15:0] _T_8465; // @[Mux.scala 31:69:@4741.4]
  wire [15:0] _T_8466; // @[Mux.scala 31:69:@4742.4]
  wire [15:0] _T_8467; // @[Mux.scala 31:69:@4743.4]
  wire [15:0] _T_8468; // @[Mux.scala 31:69:@4744.4]
  wire [15:0] _T_8469; // @[Mux.scala 31:69:@4745.4]
  wire [15:0] _T_8470; // @[Mux.scala 31:69:@4746.4]
  wire [15:0] _T_8471; // @[Mux.scala 31:69:@4747.4]
  wire [15:0] _T_8472; // @[Mux.scala 31:69:@4748.4]
  wire [15:0] _T_8473; // @[Mux.scala 31:69:@4749.4]
  wire [15:0] _T_8474; // @[Mux.scala 31:69:@4750.4]
  wire [15:0] _T_8475; // @[Mux.scala 31:69:@4751.4]
  wire [15:0] _T_8476; // @[Mux.scala 31:69:@4752.4]
  wire [15:0] _T_8477; // @[Mux.scala 31:69:@4753.4]
  wire [15:0] _T_8478; // @[Mux.scala 31:69:@4754.4]
  wire [15:0] _T_8479; // @[Mux.scala 31:69:@4755.4]
  wire [15:0] _T_8480; // @[Mux.scala 31:69:@4756.4]
  wire  _T_8481; // @[OneHot.scala 66:30:@4757.4]
  wire  _T_8482; // @[OneHot.scala 66:30:@4758.4]
  wire  _T_8483; // @[OneHot.scala 66:30:@4759.4]
  wire  _T_8484; // @[OneHot.scala 66:30:@4760.4]
  wire  _T_8485; // @[OneHot.scala 66:30:@4761.4]
  wire  _T_8486; // @[OneHot.scala 66:30:@4762.4]
  wire  _T_8487; // @[OneHot.scala 66:30:@4763.4]
  wire  _T_8488; // @[OneHot.scala 66:30:@4764.4]
  wire  _T_8489; // @[OneHot.scala 66:30:@4765.4]
  wire  _T_8490; // @[OneHot.scala 66:30:@4766.4]
  wire  _T_8491; // @[OneHot.scala 66:30:@4767.4]
  wire  _T_8492; // @[OneHot.scala 66:30:@4768.4]
  wire  _T_8493; // @[OneHot.scala 66:30:@4769.4]
  wire  _T_8494; // @[OneHot.scala 66:30:@4770.4]
  wire  _T_8495; // @[OneHot.scala 66:30:@4771.4]
  wire  _T_8496; // @[OneHot.scala 66:30:@4772.4]
  wire [15:0] _T_8537; // @[Mux.scala 31:69:@4790.4]
  wire [15:0] _T_8538; // @[Mux.scala 31:69:@4791.4]
  wire [15:0] _T_8539; // @[Mux.scala 31:69:@4792.4]
  wire [15:0] _T_8540; // @[Mux.scala 31:69:@4793.4]
  wire [15:0] _T_8541; // @[Mux.scala 31:69:@4794.4]
  wire [15:0] _T_8542; // @[Mux.scala 31:69:@4795.4]
  wire [15:0] _T_8543; // @[Mux.scala 31:69:@4796.4]
  wire [15:0] _T_8544; // @[Mux.scala 31:69:@4797.4]
  wire [15:0] _T_8545; // @[Mux.scala 31:69:@4798.4]
  wire [15:0] _T_8546; // @[Mux.scala 31:69:@4799.4]
  wire [15:0] _T_8547; // @[Mux.scala 31:69:@4800.4]
  wire [15:0] _T_8548; // @[Mux.scala 31:69:@4801.4]
  wire [15:0] _T_8549; // @[Mux.scala 31:69:@4802.4]
  wire [15:0] _T_8550; // @[Mux.scala 31:69:@4803.4]
  wire [15:0] _T_8551; // @[Mux.scala 31:69:@4804.4]
  wire [15:0] _T_8552; // @[Mux.scala 31:69:@4805.4]
  wire  _T_8553; // @[OneHot.scala 66:30:@4806.4]
  wire  _T_8554; // @[OneHot.scala 66:30:@4807.4]
  wire  _T_8555; // @[OneHot.scala 66:30:@4808.4]
  wire  _T_8556; // @[OneHot.scala 66:30:@4809.4]
  wire  _T_8557; // @[OneHot.scala 66:30:@4810.4]
  wire  _T_8558; // @[OneHot.scala 66:30:@4811.4]
  wire  _T_8559; // @[OneHot.scala 66:30:@4812.4]
  wire  _T_8560; // @[OneHot.scala 66:30:@4813.4]
  wire  _T_8561; // @[OneHot.scala 66:30:@4814.4]
  wire  _T_8562; // @[OneHot.scala 66:30:@4815.4]
  wire  _T_8563; // @[OneHot.scala 66:30:@4816.4]
  wire  _T_8564; // @[OneHot.scala 66:30:@4817.4]
  wire  _T_8565; // @[OneHot.scala 66:30:@4818.4]
  wire  _T_8566; // @[OneHot.scala 66:30:@4819.4]
  wire  _T_8567; // @[OneHot.scala 66:30:@4820.4]
  wire  _T_8568; // @[OneHot.scala 66:30:@4821.4]
  wire [15:0] _T_8609; // @[Mux.scala 31:69:@4839.4]
  wire [15:0] _T_8610; // @[Mux.scala 31:69:@4840.4]
  wire [15:0] _T_8611; // @[Mux.scala 31:69:@4841.4]
  wire [15:0] _T_8612; // @[Mux.scala 31:69:@4842.4]
  wire [15:0] _T_8613; // @[Mux.scala 31:69:@4843.4]
  wire [15:0] _T_8614; // @[Mux.scala 31:69:@4844.4]
  wire [15:0] _T_8615; // @[Mux.scala 31:69:@4845.4]
  wire [15:0] _T_8616; // @[Mux.scala 31:69:@4846.4]
  wire [15:0] _T_8617; // @[Mux.scala 31:69:@4847.4]
  wire [15:0] _T_8618; // @[Mux.scala 31:69:@4848.4]
  wire [15:0] _T_8619; // @[Mux.scala 31:69:@4849.4]
  wire [15:0] _T_8620; // @[Mux.scala 31:69:@4850.4]
  wire [15:0] _T_8621; // @[Mux.scala 31:69:@4851.4]
  wire [15:0] _T_8622; // @[Mux.scala 31:69:@4852.4]
  wire [15:0] _T_8623; // @[Mux.scala 31:69:@4853.4]
  wire [15:0] _T_8624; // @[Mux.scala 31:69:@4854.4]
  wire  _T_8625; // @[OneHot.scala 66:30:@4855.4]
  wire  _T_8626; // @[OneHot.scala 66:30:@4856.4]
  wire  _T_8627; // @[OneHot.scala 66:30:@4857.4]
  wire  _T_8628; // @[OneHot.scala 66:30:@4858.4]
  wire  _T_8629; // @[OneHot.scala 66:30:@4859.4]
  wire  _T_8630; // @[OneHot.scala 66:30:@4860.4]
  wire  _T_8631; // @[OneHot.scala 66:30:@4861.4]
  wire  _T_8632; // @[OneHot.scala 66:30:@4862.4]
  wire  _T_8633; // @[OneHot.scala 66:30:@4863.4]
  wire  _T_8634; // @[OneHot.scala 66:30:@4864.4]
  wire  _T_8635; // @[OneHot.scala 66:30:@4865.4]
  wire  _T_8636; // @[OneHot.scala 66:30:@4866.4]
  wire  _T_8637; // @[OneHot.scala 66:30:@4867.4]
  wire  _T_8638; // @[OneHot.scala 66:30:@4868.4]
  wire  _T_8639; // @[OneHot.scala 66:30:@4869.4]
  wire  _T_8640; // @[OneHot.scala 66:30:@4870.4]
  wire [15:0] _T_8681; // @[Mux.scala 31:69:@4888.4]
  wire [15:0] _T_8682; // @[Mux.scala 31:69:@4889.4]
  wire [15:0] _T_8683; // @[Mux.scala 31:69:@4890.4]
  wire [15:0] _T_8684; // @[Mux.scala 31:69:@4891.4]
  wire [15:0] _T_8685; // @[Mux.scala 31:69:@4892.4]
  wire [15:0] _T_8686; // @[Mux.scala 31:69:@4893.4]
  wire [15:0] _T_8687; // @[Mux.scala 31:69:@4894.4]
  wire [15:0] _T_8688; // @[Mux.scala 31:69:@4895.4]
  wire [15:0] _T_8689; // @[Mux.scala 31:69:@4896.4]
  wire [15:0] _T_8690; // @[Mux.scala 31:69:@4897.4]
  wire [15:0] _T_8691; // @[Mux.scala 31:69:@4898.4]
  wire [15:0] _T_8692; // @[Mux.scala 31:69:@4899.4]
  wire [15:0] _T_8693; // @[Mux.scala 31:69:@4900.4]
  wire [15:0] _T_8694; // @[Mux.scala 31:69:@4901.4]
  wire [15:0] _T_8695; // @[Mux.scala 31:69:@4902.4]
  wire [15:0] _T_8696; // @[Mux.scala 31:69:@4903.4]
  wire  _T_8697; // @[OneHot.scala 66:30:@4904.4]
  wire  _T_8698; // @[OneHot.scala 66:30:@4905.4]
  wire  _T_8699; // @[OneHot.scala 66:30:@4906.4]
  wire  _T_8700; // @[OneHot.scala 66:30:@4907.4]
  wire  _T_8701; // @[OneHot.scala 66:30:@4908.4]
  wire  _T_8702; // @[OneHot.scala 66:30:@4909.4]
  wire  _T_8703; // @[OneHot.scala 66:30:@4910.4]
  wire  _T_8704; // @[OneHot.scala 66:30:@4911.4]
  wire  _T_8705; // @[OneHot.scala 66:30:@4912.4]
  wire  _T_8706; // @[OneHot.scala 66:30:@4913.4]
  wire  _T_8707; // @[OneHot.scala 66:30:@4914.4]
  wire  _T_8708; // @[OneHot.scala 66:30:@4915.4]
  wire  _T_8709; // @[OneHot.scala 66:30:@4916.4]
  wire  _T_8710; // @[OneHot.scala 66:30:@4917.4]
  wire  _T_8711; // @[OneHot.scala 66:30:@4918.4]
  wire  _T_8712; // @[OneHot.scala 66:30:@4919.4]
  wire [15:0] _T_8753; // @[Mux.scala 31:69:@4937.4]
  wire [15:0] _T_8754; // @[Mux.scala 31:69:@4938.4]
  wire [15:0] _T_8755; // @[Mux.scala 31:69:@4939.4]
  wire [15:0] _T_8756; // @[Mux.scala 31:69:@4940.4]
  wire [15:0] _T_8757; // @[Mux.scala 31:69:@4941.4]
  wire [15:0] _T_8758; // @[Mux.scala 31:69:@4942.4]
  wire [15:0] _T_8759; // @[Mux.scala 31:69:@4943.4]
  wire [15:0] _T_8760; // @[Mux.scala 31:69:@4944.4]
  wire [15:0] _T_8761; // @[Mux.scala 31:69:@4945.4]
  wire [15:0] _T_8762; // @[Mux.scala 31:69:@4946.4]
  wire [15:0] _T_8763; // @[Mux.scala 31:69:@4947.4]
  wire [15:0] _T_8764; // @[Mux.scala 31:69:@4948.4]
  wire [15:0] _T_8765; // @[Mux.scala 31:69:@4949.4]
  wire [15:0] _T_8766; // @[Mux.scala 31:69:@4950.4]
  wire [15:0] _T_8767; // @[Mux.scala 31:69:@4951.4]
  wire [15:0] _T_8768; // @[Mux.scala 31:69:@4952.4]
  wire  _T_8769; // @[OneHot.scala 66:30:@4953.4]
  wire  _T_8770; // @[OneHot.scala 66:30:@4954.4]
  wire  _T_8771; // @[OneHot.scala 66:30:@4955.4]
  wire  _T_8772; // @[OneHot.scala 66:30:@4956.4]
  wire  _T_8773; // @[OneHot.scala 66:30:@4957.4]
  wire  _T_8774; // @[OneHot.scala 66:30:@4958.4]
  wire  _T_8775; // @[OneHot.scala 66:30:@4959.4]
  wire  _T_8776; // @[OneHot.scala 66:30:@4960.4]
  wire  _T_8777; // @[OneHot.scala 66:30:@4961.4]
  wire  _T_8778; // @[OneHot.scala 66:30:@4962.4]
  wire  _T_8779; // @[OneHot.scala 66:30:@4963.4]
  wire  _T_8780; // @[OneHot.scala 66:30:@4964.4]
  wire  _T_8781; // @[OneHot.scala 66:30:@4965.4]
  wire  _T_8782; // @[OneHot.scala 66:30:@4966.4]
  wire  _T_8783; // @[OneHot.scala 66:30:@4967.4]
  wire  _T_8784; // @[OneHot.scala 66:30:@4968.4]
  wire [15:0] _T_8825; // @[Mux.scala 31:69:@4986.4]
  wire [15:0] _T_8826; // @[Mux.scala 31:69:@4987.4]
  wire [15:0] _T_8827; // @[Mux.scala 31:69:@4988.4]
  wire [15:0] _T_8828; // @[Mux.scala 31:69:@4989.4]
  wire [15:0] _T_8829; // @[Mux.scala 31:69:@4990.4]
  wire [15:0] _T_8830; // @[Mux.scala 31:69:@4991.4]
  wire [15:0] _T_8831; // @[Mux.scala 31:69:@4992.4]
  wire [15:0] _T_8832; // @[Mux.scala 31:69:@4993.4]
  wire [15:0] _T_8833; // @[Mux.scala 31:69:@4994.4]
  wire [15:0] _T_8834; // @[Mux.scala 31:69:@4995.4]
  wire [15:0] _T_8835; // @[Mux.scala 31:69:@4996.4]
  wire [15:0] _T_8836; // @[Mux.scala 31:69:@4997.4]
  wire [15:0] _T_8837; // @[Mux.scala 31:69:@4998.4]
  wire [15:0] _T_8838; // @[Mux.scala 31:69:@4999.4]
  wire [15:0] _T_8839; // @[Mux.scala 31:69:@5000.4]
  wire [15:0] _T_8840; // @[Mux.scala 31:69:@5001.4]
  wire  _T_8841; // @[OneHot.scala 66:30:@5002.4]
  wire  _T_8842; // @[OneHot.scala 66:30:@5003.4]
  wire  _T_8843; // @[OneHot.scala 66:30:@5004.4]
  wire  _T_8844; // @[OneHot.scala 66:30:@5005.4]
  wire  _T_8845; // @[OneHot.scala 66:30:@5006.4]
  wire  _T_8846; // @[OneHot.scala 66:30:@5007.4]
  wire  _T_8847; // @[OneHot.scala 66:30:@5008.4]
  wire  _T_8848; // @[OneHot.scala 66:30:@5009.4]
  wire  _T_8849; // @[OneHot.scala 66:30:@5010.4]
  wire  _T_8850; // @[OneHot.scala 66:30:@5011.4]
  wire  _T_8851; // @[OneHot.scala 66:30:@5012.4]
  wire  _T_8852; // @[OneHot.scala 66:30:@5013.4]
  wire  _T_8853; // @[OneHot.scala 66:30:@5014.4]
  wire  _T_8854; // @[OneHot.scala 66:30:@5015.4]
  wire  _T_8855; // @[OneHot.scala 66:30:@5016.4]
  wire  _T_8856; // @[OneHot.scala 66:30:@5017.4]
  wire [15:0] _T_8897; // @[Mux.scala 31:69:@5035.4]
  wire [15:0] _T_8898; // @[Mux.scala 31:69:@5036.4]
  wire [15:0] _T_8899; // @[Mux.scala 31:69:@5037.4]
  wire [15:0] _T_8900; // @[Mux.scala 31:69:@5038.4]
  wire [15:0] _T_8901; // @[Mux.scala 31:69:@5039.4]
  wire [15:0] _T_8902; // @[Mux.scala 31:69:@5040.4]
  wire [15:0] _T_8903; // @[Mux.scala 31:69:@5041.4]
  wire [15:0] _T_8904; // @[Mux.scala 31:69:@5042.4]
  wire [15:0] _T_8905; // @[Mux.scala 31:69:@5043.4]
  wire [15:0] _T_8906; // @[Mux.scala 31:69:@5044.4]
  wire [15:0] _T_8907; // @[Mux.scala 31:69:@5045.4]
  wire [15:0] _T_8908; // @[Mux.scala 31:69:@5046.4]
  wire [15:0] _T_8909; // @[Mux.scala 31:69:@5047.4]
  wire [15:0] _T_8910; // @[Mux.scala 31:69:@5048.4]
  wire [15:0] _T_8911; // @[Mux.scala 31:69:@5049.4]
  wire [15:0] _T_8912; // @[Mux.scala 31:69:@5050.4]
  wire  _T_8913; // @[OneHot.scala 66:30:@5051.4]
  wire  _T_8914; // @[OneHot.scala 66:30:@5052.4]
  wire  _T_8915; // @[OneHot.scala 66:30:@5053.4]
  wire  _T_8916; // @[OneHot.scala 66:30:@5054.4]
  wire  _T_8917; // @[OneHot.scala 66:30:@5055.4]
  wire  _T_8918; // @[OneHot.scala 66:30:@5056.4]
  wire  _T_8919; // @[OneHot.scala 66:30:@5057.4]
  wire  _T_8920; // @[OneHot.scala 66:30:@5058.4]
  wire  _T_8921; // @[OneHot.scala 66:30:@5059.4]
  wire  _T_8922; // @[OneHot.scala 66:30:@5060.4]
  wire  _T_8923; // @[OneHot.scala 66:30:@5061.4]
  wire  _T_8924; // @[OneHot.scala 66:30:@5062.4]
  wire  _T_8925; // @[OneHot.scala 66:30:@5063.4]
  wire  _T_8926; // @[OneHot.scala 66:30:@5064.4]
  wire  _T_8927; // @[OneHot.scala 66:30:@5065.4]
  wire  _T_8928; // @[OneHot.scala 66:30:@5066.4]
  wire [15:0] _T_8969; // @[Mux.scala 31:69:@5084.4]
  wire [15:0] _T_8970; // @[Mux.scala 31:69:@5085.4]
  wire [15:0] _T_8971; // @[Mux.scala 31:69:@5086.4]
  wire [15:0] _T_8972; // @[Mux.scala 31:69:@5087.4]
  wire [15:0] _T_8973; // @[Mux.scala 31:69:@5088.4]
  wire [15:0] _T_8974; // @[Mux.scala 31:69:@5089.4]
  wire [15:0] _T_8975; // @[Mux.scala 31:69:@5090.4]
  wire [15:0] _T_8976; // @[Mux.scala 31:69:@5091.4]
  wire [15:0] _T_8977; // @[Mux.scala 31:69:@5092.4]
  wire [15:0] _T_8978; // @[Mux.scala 31:69:@5093.4]
  wire [15:0] _T_8979; // @[Mux.scala 31:69:@5094.4]
  wire [15:0] _T_8980; // @[Mux.scala 31:69:@5095.4]
  wire [15:0] _T_8981; // @[Mux.scala 31:69:@5096.4]
  wire [15:0] _T_8982; // @[Mux.scala 31:69:@5097.4]
  wire [15:0] _T_8983; // @[Mux.scala 31:69:@5098.4]
  wire [15:0] _T_8984; // @[Mux.scala 31:69:@5099.4]
  wire  _T_8985; // @[OneHot.scala 66:30:@5100.4]
  wire  _T_8986; // @[OneHot.scala 66:30:@5101.4]
  wire  _T_8987; // @[OneHot.scala 66:30:@5102.4]
  wire  _T_8988; // @[OneHot.scala 66:30:@5103.4]
  wire  _T_8989; // @[OneHot.scala 66:30:@5104.4]
  wire  _T_8990; // @[OneHot.scala 66:30:@5105.4]
  wire  _T_8991; // @[OneHot.scala 66:30:@5106.4]
  wire  _T_8992; // @[OneHot.scala 66:30:@5107.4]
  wire  _T_8993; // @[OneHot.scala 66:30:@5108.4]
  wire  _T_8994; // @[OneHot.scala 66:30:@5109.4]
  wire  _T_8995; // @[OneHot.scala 66:30:@5110.4]
  wire  _T_8996; // @[OneHot.scala 66:30:@5111.4]
  wire  _T_8997; // @[OneHot.scala 66:30:@5112.4]
  wire  _T_8998; // @[OneHot.scala 66:30:@5113.4]
  wire  _T_8999; // @[OneHot.scala 66:30:@5114.4]
  wire  _T_9000; // @[OneHot.scala 66:30:@5115.4]
  wire [15:0] _T_9041; // @[Mux.scala 31:69:@5133.4]
  wire [15:0] _T_9042; // @[Mux.scala 31:69:@5134.4]
  wire [15:0] _T_9043; // @[Mux.scala 31:69:@5135.4]
  wire [15:0] _T_9044; // @[Mux.scala 31:69:@5136.4]
  wire [15:0] _T_9045; // @[Mux.scala 31:69:@5137.4]
  wire [15:0] _T_9046; // @[Mux.scala 31:69:@5138.4]
  wire [15:0] _T_9047; // @[Mux.scala 31:69:@5139.4]
  wire [15:0] _T_9048; // @[Mux.scala 31:69:@5140.4]
  wire [15:0] _T_9049; // @[Mux.scala 31:69:@5141.4]
  wire [15:0] _T_9050; // @[Mux.scala 31:69:@5142.4]
  wire [15:0] _T_9051; // @[Mux.scala 31:69:@5143.4]
  wire [15:0] _T_9052; // @[Mux.scala 31:69:@5144.4]
  wire [15:0] _T_9053; // @[Mux.scala 31:69:@5145.4]
  wire [15:0] _T_9054; // @[Mux.scala 31:69:@5146.4]
  wire [15:0] _T_9055; // @[Mux.scala 31:69:@5147.4]
  wire [15:0] _T_9056; // @[Mux.scala 31:69:@5148.4]
  wire  _T_9057; // @[OneHot.scala 66:30:@5149.4]
  wire  _T_9058; // @[OneHot.scala 66:30:@5150.4]
  wire  _T_9059; // @[OneHot.scala 66:30:@5151.4]
  wire  _T_9060; // @[OneHot.scala 66:30:@5152.4]
  wire  _T_9061; // @[OneHot.scala 66:30:@5153.4]
  wire  _T_9062; // @[OneHot.scala 66:30:@5154.4]
  wire  _T_9063; // @[OneHot.scala 66:30:@5155.4]
  wire  _T_9064; // @[OneHot.scala 66:30:@5156.4]
  wire  _T_9065; // @[OneHot.scala 66:30:@5157.4]
  wire  _T_9066; // @[OneHot.scala 66:30:@5158.4]
  wire  _T_9067; // @[OneHot.scala 66:30:@5159.4]
  wire  _T_9068; // @[OneHot.scala 66:30:@5160.4]
  wire  _T_9069; // @[OneHot.scala 66:30:@5161.4]
  wire  _T_9070; // @[OneHot.scala 66:30:@5162.4]
  wire  _T_9071; // @[OneHot.scala 66:30:@5163.4]
  wire  _T_9072; // @[OneHot.scala 66:30:@5164.4]
  wire [15:0] _T_9113; // @[Mux.scala 31:69:@5182.4]
  wire [15:0] _T_9114; // @[Mux.scala 31:69:@5183.4]
  wire [15:0] _T_9115; // @[Mux.scala 31:69:@5184.4]
  wire [15:0] _T_9116; // @[Mux.scala 31:69:@5185.4]
  wire [15:0] _T_9117; // @[Mux.scala 31:69:@5186.4]
  wire [15:0] _T_9118; // @[Mux.scala 31:69:@5187.4]
  wire [15:0] _T_9119; // @[Mux.scala 31:69:@5188.4]
  wire [15:0] _T_9120; // @[Mux.scala 31:69:@5189.4]
  wire [15:0] _T_9121; // @[Mux.scala 31:69:@5190.4]
  wire [15:0] _T_9122; // @[Mux.scala 31:69:@5191.4]
  wire [15:0] _T_9123; // @[Mux.scala 31:69:@5192.4]
  wire [15:0] _T_9124; // @[Mux.scala 31:69:@5193.4]
  wire [15:0] _T_9125; // @[Mux.scala 31:69:@5194.4]
  wire [15:0] _T_9126; // @[Mux.scala 31:69:@5195.4]
  wire [15:0] _T_9127; // @[Mux.scala 31:69:@5196.4]
  wire [15:0] _T_9128; // @[Mux.scala 31:69:@5197.4]
  wire  _T_9129; // @[OneHot.scala 66:30:@5198.4]
  wire  _T_9130; // @[OneHot.scala 66:30:@5199.4]
  wire  _T_9131; // @[OneHot.scala 66:30:@5200.4]
  wire  _T_9132; // @[OneHot.scala 66:30:@5201.4]
  wire  _T_9133; // @[OneHot.scala 66:30:@5202.4]
  wire  _T_9134; // @[OneHot.scala 66:30:@5203.4]
  wire  _T_9135; // @[OneHot.scala 66:30:@5204.4]
  wire  _T_9136; // @[OneHot.scala 66:30:@5205.4]
  wire  _T_9137; // @[OneHot.scala 66:30:@5206.4]
  wire  _T_9138; // @[OneHot.scala 66:30:@5207.4]
  wire  _T_9139; // @[OneHot.scala 66:30:@5208.4]
  wire  _T_9140; // @[OneHot.scala 66:30:@5209.4]
  wire  _T_9141; // @[OneHot.scala 66:30:@5210.4]
  wire  _T_9142; // @[OneHot.scala 66:30:@5211.4]
  wire  _T_9143; // @[OneHot.scala 66:30:@5212.4]
  wire  _T_9144; // @[OneHot.scala 66:30:@5213.4]
  wire [7:0] _T_9209; // @[Mux.scala 19:72:@5237.4]
  wire [15:0] _T_9217; // @[Mux.scala 19:72:@5245.4]
  wire [15:0] _T_9219; // @[Mux.scala 19:72:@5246.4]
  wire [7:0] _T_9226; // @[Mux.scala 19:72:@5253.4]
  wire [15:0] _T_9234; // @[Mux.scala 19:72:@5261.4]
  wire [15:0] _T_9236; // @[Mux.scala 19:72:@5262.4]
  wire [7:0] _T_9243; // @[Mux.scala 19:72:@5269.4]
  wire [15:0] _T_9251; // @[Mux.scala 19:72:@5277.4]
  wire [15:0] _T_9253; // @[Mux.scala 19:72:@5278.4]
  wire [7:0] _T_9260; // @[Mux.scala 19:72:@5285.4]
  wire [15:0] _T_9268; // @[Mux.scala 19:72:@5293.4]
  wire [15:0] _T_9270; // @[Mux.scala 19:72:@5294.4]
  wire [7:0] _T_9277; // @[Mux.scala 19:72:@5301.4]
  wire [15:0] _T_9285; // @[Mux.scala 19:72:@5309.4]
  wire [15:0] _T_9287; // @[Mux.scala 19:72:@5310.4]
  wire [7:0] _T_9294; // @[Mux.scala 19:72:@5317.4]
  wire [15:0] _T_9302; // @[Mux.scala 19:72:@5325.4]
  wire [15:0] _T_9304; // @[Mux.scala 19:72:@5326.4]
  wire [7:0] _T_9311; // @[Mux.scala 19:72:@5333.4]
  wire [15:0] _T_9319; // @[Mux.scala 19:72:@5341.4]
  wire [15:0] _T_9321; // @[Mux.scala 19:72:@5342.4]
  wire [7:0] _T_9328; // @[Mux.scala 19:72:@5349.4]
  wire [15:0] _T_9336; // @[Mux.scala 19:72:@5357.4]
  wire [15:0] _T_9338; // @[Mux.scala 19:72:@5358.4]
  wire [7:0] _T_9345; // @[Mux.scala 19:72:@5365.4]
  wire [15:0] _T_9353; // @[Mux.scala 19:72:@5373.4]
  wire [15:0] _T_9355; // @[Mux.scala 19:72:@5374.4]
  wire [7:0] _T_9362; // @[Mux.scala 19:72:@5381.4]
  wire [15:0] _T_9370; // @[Mux.scala 19:72:@5389.4]
  wire [15:0] _T_9372; // @[Mux.scala 19:72:@5390.4]
  wire [7:0] _T_9379; // @[Mux.scala 19:72:@5397.4]
  wire [15:0] _T_9387; // @[Mux.scala 19:72:@5405.4]
  wire [15:0] _T_9389; // @[Mux.scala 19:72:@5406.4]
  wire [7:0] _T_9396; // @[Mux.scala 19:72:@5413.4]
  wire [15:0] _T_9404; // @[Mux.scala 19:72:@5421.4]
  wire [15:0] _T_9406; // @[Mux.scala 19:72:@5422.4]
  wire [7:0] _T_9413; // @[Mux.scala 19:72:@5429.4]
  wire [15:0] _T_9421; // @[Mux.scala 19:72:@5437.4]
  wire [15:0] _T_9423; // @[Mux.scala 19:72:@5438.4]
  wire [7:0] _T_9430; // @[Mux.scala 19:72:@5445.4]
  wire [15:0] _T_9438; // @[Mux.scala 19:72:@5453.4]
  wire [15:0] _T_9440; // @[Mux.scala 19:72:@5454.4]
  wire [7:0] _T_9447; // @[Mux.scala 19:72:@5461.4]
  wire [15:0] _T_9455; // @[Mux.scala 19:72:@5469.4]
  wire [15:0] _T_9457; // @[Mux.scala 19:72:@5470.4]
  wire [7:0] _T_9464; // @[Mux.scala 19:72:@5477.4]
  wire [15:0] _T_9472; // @[Mux.scala 19:72:@5485.4]
  wire [15:0] _T_9474; // @[Mux.scala 19:72:@5486.4]
  wire [15:0] _T_9475; // @[Mux.scala 19:72:@5487.4]
  wire [15:0] _T_9476; // @[Mux.scala 19:72:@5488.4]
  wire [15:0] _T_9477; // @[Mux.scala 19:72:@5489.4]
  wire [15:0] _T_9478; // @[Mux.scala 19:72:@5490.4]
  wire [15:0] _T_9479; // @[Mux.scala 19:72:@5491.4]
  wire [15:0] _T_9480; // @[Mux.scala 19:72:@5492.4]
  wire [15:0] _T_9481; // @[Mux.scala 19:72:@5493.4]
  wire [15:0] _T_9482; // @[Mux.scala 19:72:@5494.4]
  wire [15:0] _T_9483; // @[Mux.scala 19:72:@5495.4]
  wire [15:0] _T_9484; // @[Mux.scala 19:72:@5496.4]
  wire [15:0] _T_9485; // @[Mux.scala 19:72:@5497.4]
  wire [15:0] _T_9486; // @[Mux.scala 19:72:@5498.4]
  wire [15:0] _T_9487; // @[Mux.scala 19:72:@5499.4]
  wire [15:0] _T_9488; // @[Mux.scala 19:72:@5500.4]
  wire [15:0] _T_9489; // @[Mux.scala 19:72:@5501.4]
  wire  inputAddrPriorityPorts_1_0; // @[Mux.scala 19:72:@5505.4]
  wire  inputAddrPriorityPorts_1_1; // @[Mux.scala 19:72:@5507.4]
  wire  inputAddrPriorityPorts_1_2; // @[Mux.scala 19:72:@5509.4]
  wire  inputAddrPriorityPorts_1_3; // @[Mux.scala 19:72:@5511.4]
  wire  inputAddrPriorityPorts_1_4; // @[Mux.scala 19:72:@5513.4]
  wire  inputAddrPriorityPorts_1_5; // @[Mux.scala 19:72:@5515.4]
  wire  inputAddrPriorityPorts_1_6; // @[Mux.scala 19:72:@5517.4]
  wire  inputAddrPriorityPorts_1_7; // @[Mux.scala 19:72:@5519.4]
  wire  inputAddrPriorityPorts_1_8; // @[Mux.scala 19:72:@5521.4]
  wire  inputAddrPriorityPorts_1_9; // @[Mux.scala 19:72:@5523.4]
  wire  inputAddrPriorityPorts_1_10; // @[Mux.scala 19:72:@5525.4]
  wire  inputAddrPriorityPorts_1_11; // @[Mux.scala 19:72:@5527.4]
  wire  inputAddrPriorityPorts_1_12; // @[Mux.scala 19:72:@5529.4]
  wire  inputAddrPriorityPorts_1_13; // @[Mux.scala 19:72:@5531.4]
  wire  inputAddrPriorityPorts_1_14; // @[Mux.scala 19:72:@5533.4]
  wire  inputAddrPriorityPorts_1_15; // @[Mux.scala 19:72:@5535.4]
  wire [15:0] _T_9691; // @[Mux.scala 31:69:@5589.4]
  wire [15:0] _T_9692; // @[Mux.scala 31:69:@5590.4]
  wire [15:0] _T_9693; // @[Mux.scala 31:69:@5591.4]
  wire [15:0] _T_9694; // @[Mux.scala 31:69:@5592.4]
  wire [15:0] _T_9695; // @[Mux.scala 31:69:@5593.4]
  wire [15:0] _T_9696; // @[Mux.scala 31:69:@5594.4]
  wire [15:0] _T_9697; // @[Mux.scala 31:69:@5595.4]
  wire [15:0] _T_9698; // @[Mux.scala 31:69:@5596.4]
  wire [15:0] _T_9699; // @[Mux.scala 31:69:@5597.4]
  wire [15:0] _T_9700; // @[Mux.scala 31:69:@5598.4]
  wire [15:0] _T_9701; // @[Mux.scala 31:69:@5599.4]
  wire [15:0] _T_9702; // @[Mux.scala 31:69:@5600.4]
  wire [15:0] _T_9703; // @[Mux.scala 31:69:@5601.4]
  wire [15:0] _T_9704; // @[Mux.scala 31:69:@5602.4]
  wire [15:0] _T_9705; // @[Mux.scala 31:69:@5603.4]
  wire [15:0] _T_9706; // @[Mux.scala 31:69:@5604.4]
  wire  _T_9707; // @[OneHot.scala 66:30:@5605.4]
  wire  _T_9708; // @[OneHot.scala 66:30:@5606.4]
  wire  _T_9709; // @[OneHot.scala 66:30:@5607.4]
  wire  _T_9710; // @[OneHot.scala 66:30:@5608.4]
  wire  _T_9711; // @[OneHot.scala 66:30:@5609.4]
  wire  _T_9712; // @[OneHot.scala 66:30:@5610.4]
  wire  _T_9713; // @[OneHot.scala 66:30:@5611.4]
  wire  _T_9714; // @[OneHot.scala 66:30:@5612.4]
  wire  _T_9715; // @[OneHot.scala 66:30:@5613.4]
  wire  _T_9716; // @[OneHot.scala 66:30:@5614.4]
  wire  _T_9717; // @[OneHot.scala 66:30:@5615.4]
  wire  _T_9718; // @[OneHot.scala 66:30:@5616.4]
  wire  _T_9719; // @[OneHot.scala 66:30:@5617.4]
  wire  _T_9720; // @[OneHot.scala 66:30:@5618.4]
  wire  _T_9721; // @[OneHot.scala 66:30:@5619.4]
  wire  _T_9722; // @[OneHot.scala 66:30:@5620.4]
  wire [15:0] _T_9763; // @[Mux.scala 31:69:@5638.4]
  wire [15:0] _T_9764; // @[Mux.scala 31:69:@5639.4]
  wire [15:0] _T_9765; // @[Mux.scala 31:69:@5640.4]
  wire [15:0] _T_9766; // @[Mux.scala 31:69:@5641.4]
  wire [15:0] _T_9767; // @[Mux.scala 31:69:@5642.4]
  wire [15:0] _T_9768; // @[Mux.scala 31:69:@5643.4]
  wire [15:0] _T_9769; // @[Mux.scala 31:69:@5644.4]
  wire [15:0] _T_9770; // @[Mux.scala 31:69:@5645.4]
  wire [15:0] _T_9771; // @[Mux.scala 31:69:@5646.4]
  wire [15:0] _T_9772; // @[Mux.scala 31:69:@5647.4]
  wire [15:0] _T_9773; // @[Mux.scala 31:69:@5648.4]
  wire [15:0] _T_9774; // @[Mux.scala 31:69:@5649.4]
  wire [15:0] _T_9775; // @[Mux.scala 31:69:@5650.4]
  wire [15:0] _T_9776; // @[Mux.scala 31:69:@5651.4]
  wire [15:0] _T_9777; // @[Mux.scala 31:69:@5652.4]
  wire [15:0] _T_9778; // @[Mux.scala 31:69:@5653.4]
  wire  _T_9779; // @[OneHot.scala 66:30:@5654.4]
  wire  _T_9780; // @[OneHot.scala 66:30:@5655.4]
  wire  _T_9781; // @[OneHot.scala 66:30:@5656.4]
  wire  _T_9782; // @[OneHot.scala 66:30:@5657.4]
  wire  _T_9783; // @[OneHot.scala 66:30:@5658.4]
  wire  _T_9784; // @[OneHot.scala 66:30:@5659.4]
  wire  _T_9785; // @[OneHot.scala 66:30:@5660.4]
  wire  _T_9786; // @[OneHot.scala 66:30:@5661.4]
  wire  _T_9787; // @[OneHot.scala 66:30:@5662.4]
  wire  _T_9788; // @[OneHot.scala 66:30:@5663.4]
  wire  _T_9789; // @[OneHot.scala 66:30:@5664.4]
  wire  _T_9790; // @[OneHot.scala 66:30:@5665.4]
  wire  _T_9791; // @[OneHot.scala 66:30:@5666.4]
  wire  _T_9792; // @[OneHot.scala 66:30:@5667.4]
  wire  _T_9793; // @[OneHot.scala 66:30:@5668.4]
  wire  _T_9794; // @[OneHot.scala 66:30:@5669.4]
  wire [15:0] _T_9835; // @[Mux.scala 31:69:@5687.4]
  wire [15:0] _T_9836; // @[Mux.scala 31:69:@5688.4]
  wire [15:0] _T_9837; // @[Mux.scala 31:69:@5689.4]
  wire [15:0] _T_9838; // @[Mux.scala 31:69:@5690.4]
  wire [15:0] _T_9839; // @[Mux.scala 31:69:@5691.4]
  wire [15:0] _T_9840; // @[Mux.scala 31:69:@5692.4]
  wire [15:0] _T_9841; // @[Mux.scala 31:69:@5693.4]
  wire [15:0] _T_9842; // @[Mux.scala 31:69:@5694.4]
  wire [15:0] _T_9843; // @[Mux.scala 31:69:@5695.4]
  wire [15:0] _T_9844; // @[Mux.scala 31:69:@5696.4]
  wire [15:0] _T_9845; // @[Mux.scala 31:69:@5697.4]
  wire [15:0] _T_9846; // @[Mux.scala 31:69:@5698.4]
  wire [15:0] _T_9847; // @[Mux.scala 31:69:@5699.4]
  wire [15:0] _T_9848; // @[Mux.scala 31:69:@5700.4]
  wire [15:0] _T_9849; // @[Mux.scala 31:69:@5701.4]
  wire [15:0] _T_9850; // @[Mux.scala 31:69:@5702.4]
  wire  _T_9851; // @[OneHot.scala 66:30:@5703.4]
  wire  _T_9852; // @[OneHot.scala 66:30:@5704.4]
  wire  _T_9853; // @[OneHot.scala 66:30:@5705.4]
  wire  _T_9854; // @[OneHot.scala 66:30:@5706.4]
  wire  _T_9855; // @[OneHot.scala 66:30:@5707.4]
  wire  _T_9856; // @[OneHot.scala 66:30:@5708.4]
  wire  _T_9857; // @[OneHot.scala 66:30:@5709.4]
  wire  _T_9858; // @[OneHot.scala 66:30:@5710.4]
  wire  _T_9859; // @[OneHot.scala 66:30:@5711.4]
  wire  _T_9860; // @[OneHot.scala 66:30:@5712.4]
  wire  _T_9861; // @[OneHot.scala 66:30:@5713.4]
  wire  _T_9862; // @[OneHot.scala 66:30:@5714.4]
  wire  _T_9863; // @[OneHot.scala 66:30:@5715.4]
  wire  _T_9864; // @[OneHot.scala 66:30:@5716.4]
  wire  _T_9865; // @[OneHot.scala 66:30:@5717.4]
  wire  _T_9866; // @[OneHot.scala 66:30:@5718.4]
  wire [15:0] _T_9907; // @[Mux.scala 31:69:@5736.4]
  wire [15:0] _T_9908; // @[Mux.scala 31:69:@5737.4]
  wire [15:0] _T_9909; // @[Mux.scala 31:69:@5738.4]
  wire [15:0] _T_9910; // @[Mux.scala 31:69:@5739.4]
  wire [15:0] _T_9911; // @[Mux.scala 31:69:@5740.4]
  wire [15:0] _T_9912; // @[Mux.scala 31:69:@5741.4]
  wire [15:0] _T_9913; // @[Mux.scala 31:69:@5742.4]
  wire [15:0] _T_9914; // @[Mux.scala 31:69:@5743.4]
  wire [15:0] _T_9915; // @[Mux.scala 31:69:@5744.4]
  wire [15:0] _T_9916; // @[Mux.scala 31:69:@5745.4]
  wire [15:0] _T_9917; // @[Mux.scala 31:69:@5746.4]
  wire [15:0] _T_9918; // @[Mux.scala 31:69:@5747.4]
  wire [15:0] _T_9919; // @[Mux.scala 31:69:@5748.4]
  wire [15:0] _T_9920; // @[Mux.scala 31:69:@5749.4]
  wire [15:0] _T_9921; // @[Mux.scala 31:69:@5750.4]
  wire [15:0] _T_9922; // @[Mux.scala 31:69:@5751.4]
  wire  _T_9923; // @[OneHot.scala 66:30:@5752.4]
  wire  _T_9924; // @[OneHot.scala 66:30:@5753.4]
  wire  _T_9925; // @[OneHot.scala 66:30:@5754.4]
  wire  _T_9926; // @[OneHot.scala 66:30:@5755.4]
  wire  _T_9927; // @[OneHot.scala 66:30:@5756.4]
  wire  _T_9928; // @[OneHot.scala 66:30:@5757.4]
  wire  _T_9929; // @[OneHot.scala 66:30:@5758.4]
  wire  _T_9930; // @[OneHot.scala 66:30:@5759.4]
  wire  _T_9931; // @[OneHot.scala 66:30:@5760.4]
  wire  _T_9932; // @[OneHot.scala 66:30:@5761.4]
  wire  _T_9933; // @[OneHot.scala 66:30:@5762.4]
  wire  _T_9934; // @[OneHot.scala 66:30:@5763.4]
  wire  _T_9935; // @[OneHot.scala 66:30:@5764.4]
  wire  _T_9936; // @[OneHot.scala 66:30:@5765.4]
  wire  _T_9937; // @[OneHot.scala 66:30:@5766.4]
  wire  _T_9938; // @[OneHot.scala 66:30:@5767.4]
  wire [15:0] _T_9979; // @[Mux.scala 31:69:@5785.4]
  wire [15:0] _T_9980; // @[Mux.scala 31:69:@5786.4]
  wire [15:0] _T_9981; // @[Mux.scala 31:69:@5787.4]
  wire [15:0] _T_9982; // @[Mux.scala 31:69:@5788.4]
  wire [15:0] _T_9983; // @[Mux.scala 31:69:@5789.4]
  wire [15:0] _T_9984; // @[Mux.scala 31:69:@5790.4]
  wire [15:0] _T_9985; // @[Mux.scala 31:69:@5791.4]
  wire [15:0] _T_9986; // @[Mux.scala 31:69:@5792.4]
  wire [15:0] _T_9987; // @[Mux.scala 31:69:@5793.4]
  wire [15:0] _T_9988; // @[Mux.scala 31:69:@5794.4]
  wire [15:0] _T_9989; // @[Mux.scala 31:69:@5795.4]
  wire [15:0] _T_9990; // @[Mux.scala 31:69:@5796.4]
  wire [15:0] _T_9991; // @[Mux.scala 31:69:@5797.4]
  wire [15:0] _T_9992; // @[Mux.scala 31:69:@5798.4]
  wire [15:0] _T_9993; // @[Mux.scala 31:69:@5799.4]
  wire [15:0] _T_9994; // @[Mux.scala 31:69:@5800.4]
  wire  _T_9995; // @[OneHot.scala 66:30:@5801.4]
  wire  _T_9996; // @[OneHot.scala 66:30:@5802.4]
  wire  _T_9997; // @[OneHot.scala 66:30:@5803.4]
  wire  _T_9998; // @[OneHot.scala 66:30:@5804.4]
  wire  _T_9999; // @[OneHot.scala 66:30:@5805.4]
  wire  _T_10000; // @[OneHot.scala 66:30:@5806.4]
  wire  _T_10001; // @[OneHot.scala 66:30:@5807.4]
  wire  _T_10002; // @[OneHot.scala 66:30:@5808.4]
  wire  _T_10003; // @[OneHot.scala 66:30:@5809.4]
  wire  _T_10004; // @[OneHot.scala 66:30:@5810.4]
  wire  _T_10005; // @[OneHot.scala 66:30:@5811.4]
  wire  _T_10006; // @[OneHot.scala 66:30:@5812.4]
  wire  _T_10007; // @[OneHot.scala 66:30:@5813.4]
  wire  _T_10008; // @[OneHot.scala 66:30:@5814.4]
  wire  _T_10009; // @[OneHot.scala 66:30:@5815.4]
  wire  _T_10010; // @[OneHot.scala 66:30:@5816.4]
  wire [15:0] _T_10051; // @[Mux.scala 31:69:@5834.4]
  wire [15:0] _T_10052; // @[Mux.scala 31:69:@5835.4]
  wire [15:0] _T_10053; // @[Mux.scala 31:69:@5836.4]
  wire [15:0] _T_10054; // @[Mux.scala 31:69:@5837.4]
  wire [15:0] _T_10055; // @[Mux.scala 31:69:@5838.4]
  wire [15:0] _T_10056; // @[Mux.scala 31:69:@5839.4]
  wire [15:0] _T_10057; // @[Mux.scala 31:69:@5840.4]
  wire [15:0] _T_10058; // @[Mux.scala 31:69:@5841.4]
  wire [15:0] _T_10059; // @[Mux.scala 31:69:@5842.4]
  wire [15:0] _T_10060; // @[Mux.scala 31:69:@5843.4]
  wire [15:0] _T_10061; // @[Mux.scala 31:69:@5844.4]
  wire [15:0] _T_10062; // @[Mux.scala 31:69:@5845.4]
  wire [15:0] _T_10063; // @[Mux.scala 31:69:@5846.4]
  wire [15:0] _T_10064; // @[Mux.scala 31:69:@5847.4]
  wire [15:0] _T_10065; // @[Mux.scala 31:69:@5848.4]
  wire [15:0] _T_10066; // @[Mux.scala 31:69:@5849.4]
  wire  _T_10067; // @[OneHot.scala 66:30:@5850.4]
  wire  _T_10068; // @[OneHot.scala 66:30:@5851.4]
  wire  _T_10069; // @[OneHot.scala 66:30:@5852.4]
  wire  _T_10070; // @[OneHot.scala 66:30:@5853.4]
  wire  _T_10071; // @[OneHot.scala 66:30:@5854.4]
  wire  _T_10072; // @[OneHot.scala 66:30:@5855.4]
  wire  _T_10073; // @[OneHot.scala 66:30:@5856.4]
  wire  _T_10074; // @[OneHot.scala 66:30:@5857.4]
  wire  _T_10075; // @[OneHot.scala 66:30:@5858.4]
  wire  _T_10076; // @[OneHot.scala 66:30:@5859.4]
  wire  _T_10077; // @[OneHot.scala 66:30:@5860.4]
  wire  _T_10078; // @[OneHot.scala 66:30:@5861.4]
  wire  _T_10079; // @[OneHot.scala 66:30:@5862.4]
  wire  _T_10080; // @[OneHot.scala 66:30:@5863.4]
  wire  _T_10081; // @[OneHot.scala 66:30:@5864.4]
  wire  _T_10082; // @[OneHot.scala 66:30:@5865.4]
  wire [15:0] _T_10123; // @[Mux.scala 31:69:@5883.4]
  wire [15:0] _T_10124; // @[Mux.scala 31:69:@5884.4]
  wire [15:0] _T_10125; // @[Mux.scala 31:69:@5885.4]
  wire [15:0] _T_10126; // @[Mux.scala 31:69:@5886.4]
  wire [15:0] _T_10127; // @[Mux.scala 31:69:@5887.4]
  wire [15:0] _T_10128; // @[Mux.scala 31:69:@5888.4]
  wire [15:0] _T_10129; // @[Mux.scala 31:69:@5889.4]
  wire [15:0] _T_10130; // @[Mux.scala 31:69:@5890.4]
  wire [15:0] _T_10131; // @[Mux.scala 31:69:@5891.4]
  wire [15:0] _T_10132; // @[Mux.scala 31:69:@5892.4]
  wire [15:0] _T_10133; // @[Mux.scala 31:69:@5893.4]
  wire [15:0] _T_10134; // @[Mux.scala 31:69:@5894.4]
  wire [15:0] _T_10135; // @[Mux.scala 31:69:@5895.4]
  wire [15:0] _T_10136; // @[Mux.scala 31:69:@5896.4]
  wire [15:0] _T_10137; // @[Mux.scala 31:69:@5897.4]
  wire [15:0] _T_10138; // @[Mux.scala 31:69:@5898.4]
  wire  _T_10139; // @[OneHot.scala 66:30:@5899.4]
  wire  _T_10140; // @[OneHot.scala 66:30:@5900.4]
  wire  _T_10141; // @[OneHot.scala 66:30:@5901.4]
  wire  _T_10142; // @[OneHot.scala 66:30:@5902.4]
  wire  _T_10143; // @[OneHot.scala 66:30:@5903.4]
  wire  _T_10144; // @[OneHot.scala 66:30:@5904.4]
  wire  _T_10145; // @[OneHot.scala 66:30:@5905.4]
  wire  _T_10146; // @[OneHot.scala 66:30:@5906.4]
  wire  _T_10147; // @[OneHot.scala 66:30:@5907.4]
  wire  _T_10148; // @[OneHot.scala 66:30:@5908.4]
  wire  _T_10149; // @[OneHot.scala 66:30:@5909.4]
  wire  _T_10150; // @[OneHot.scala 66:30:@5910.4]
  wire  _T_10151; // @[OneHot.scala 66:30:@5911.4]
  wire  _T_10152; // @[OneHot.scala 66:30:@5912.4]
  wire  _T_10153; // @[OneHot.scala 66:30:@5913.4]
  wire  _T_10154; // @[OneHot.scala 66:30:@5914.4]
  wire [15:0] _T_10195; // @[Mux.scala 31:69:@5932.4]
  wire [15:0] _T_10196; // @[Mux.scala 31:69:@5933.4]
  wire [15:0] _T_10197; // @[Mux.scala 31:69:@5934.4]
  wire [15:0] _T_10198; // @[Mux.scala 31:69:@5935.4]
  wire [15:0] _T_10199; // @[Mux.scala 31:69:@5936.4]
  wire [15:0] _T_10200; // @[Mux.scala 31:69:@5937.4]
  wire [15:0] _T_10201; // @[Mux.scala 31:69:@5938.4]
  wire [15:0] _T_10202; // @[Mux.scala 31:69:@5939.4]
  wire [15:0] _T_10203; // @[Mux.scala 31:69:@5940.4]
  wire [15:0] _T_10204; // @[Mux.scala 31:69:@5941.4]
  wire [15:0] _T_10205; // @[Mux.scala 31:69:@5942.4]
  wire [15:0] _T_10206; // @[Mux.scala 31:69:@5943.4]
  wire [15:0] _T_10207; // @[Mux.scala 31:69:@5944.4]
  wire [15:0] _T_10208; // @[Mux.scala 31:69:@5945.4]
  wire [15:0] _T_10209; // @[Mux.scala 31:69:@5946.4]
  wire [15:0] _T_10210; // @[Mux.scala 31:69:@5947.4]
  wire  _T_10211; // @[OneHot.scala 66:30:@5948.4]
  wire  _T_10212; // @[OneHot.scala 66:30:@5949.4]
  wire  _T_10213; // @[OneHot.scala 66:30:@5950.4]
  wire  _T_10214; // @[OneHot.scala 66:30:@5951.4]
  wire  _T_10215; // @[OneHot.scala 66:30:@5952.4]
  wire  _T_10216; // @[OneHot.scala 66:30:@5953.4]
  wire  _T_10217; // @[OneHot.scala 66:30:@5954.4]
  wire  _T_10218; // @[OneHot.scala 66:30:@5955.4]
  wire  _T_10219; // @[OneHot.scala 66:30:@5956.4]
  wire  _T_10220; // @[OneHot.scala 66:30:@5957.4]
  wire  _T_10221; // @[OneHot.scala 66:30:@5958.4]
  wire  _T_10222; // @[OneHot.scala 66:30:@5959.4]
  wire  _T_10223; // @[OneHot.scala 66:30:@5960.4]
  wire  _T_10224; // @[OneHot.scala 66:30:@5961.4]
  wire  _T_10225; // @[OneHot.scala 66:30:@5962.4]
  wire  _T_10226; // @[OneHot.scala 66:30:@5963.4]
  wire [15:0] _T_10267; // @[Mux.scala 31:69:@5981.4]
  wire [15:0] _T_10268; // @[Mux.scala 31:69:@5982.4]
  wire [15:0] _T_10269; // @[Mux.scala 31:69:@5983.4]
  wire [15:0] _T_10270; // @[Mux.scala 31:69:@5984.4]
  wire [15:0] _T_10271; // @[Mux.scala 31:69:@5985.4]
  wire [15:0] _T_10272; // @[Mux.scala 31:69:@5986.4]
  wire [15:0] _T_10273; // @[Mux.scala 31:69:@5987.4]
  wire [15:0] _T_10274; // @[Mux.scala 31:69:@5988.4]
  wire [15:0] _T_10275; // @[Mux.scala 31:69:@5989.4]
  wire [15:0] _T_10276; // @[Mux.scala 31:69:@5990.4]
  wire [15:0] _T_10277; // @[Mux.scala 31:69:@5991.4]
  wire [15:0] _T_10278; // @[Mux.scala 31:69:@5992.4]
  wire [15:0] _T_10279; // @[Mux.scala 31:69:@5993.4]
  wire [15:0] _T_10280; // @[Mux.scala 31:69:@5994.4]
  wire [15:0] _T_10281; // @[Mux.scala 31:69:@5995.4]
  wire [15:0] _T_10282; // @[Mux.scala 31:69:@5996.4]
  wire  _T_10283; // @[OneHot.scala 66:30:@5997.4]
  wire  _T_10284; // @[OneHot.scala 66:30:@5998.4]
  wire  _T_10285; // @[OneHot.scala 66:30:@5999.4]
  wire  _T_10286; // @[OneHot.scala 66:30:@6000.4]
  wire  _T_10287; // @[OneHot.scala 66:30:@6001.4]
  wire  _T_10288; // @[OneHot.scala 66:30:@6002.4]
  wire  _T_10289; // @[OneHot.scala 66:30:@6003.4]
  wire  _T_10290; // @[OneHot.scala 66:30:@6004.4]
  wire  _T_10291; // @[OneHot.scala 66:30:@6005.4]
  wire  _T_10292; // @[OneHot.scala 66:30:@6006.4]
  wire  _T_10293; // @[OneHot.scala 66:30:@6007.4]
  wire  _T_10294; // @[OneHot.scala 66:30:@6008.4]
  wire  _T_10295; // @[OneHot.scala 66:30:@6009.4]
  wire  _T_10296; // @[OneHot.scala 66:30:@6010.4]
  wire  _T_10297; // @[OneHot.scala 66:30:@6011.4]
  wire  _T_10298; // @[OneHot.scala 66:30:@6012.4]
  wire [15:0] _T_10339; // @[Mux.scala 31:69:@6030.4]
  wire [15:0] _T_10340; // @[Mux.scala 31:69:@6031.4]
  wire [15:0] _T_10341; // @[Mux.scala 31:69:@6032.4]
  wire [15:0] _T_10342; // @[Mux.scala 31:69:@6033.4]
  wire [15:0] _T_10343; // @[Mux.scala 31:69:@6034.4]
  wire [15:0] _T_10344; // @[Mux.scala 31:69:@6035.4]
  wire [15:0] _T_10345; // @[Mux.scala 31:69:@6036.4]
  wire [15:0] _T_10346; // @[Mux.scala 31:69:@6037.4]
  wire [15:0] _T_10347; // @[Mux.scala 31:69:@6038.4]
  wire [15:0] _T_10348; // @[Mux.scala 31:69:@6039.4]
  wire [15:0] _T_10349; // @[Mux.scala 31:69:@6040.4]
  wire [15:0] _T_10350; // @[Mux.scala 31:69:@6041.4]
  wire [15:0] _T_10351; // @[Mux.scala 31:69:@6042.4]
  wire [15:0] _T_10352; // @[Mux.scala 31:69:@6043.4]
  wire [15:0] _T_10353; // @[Mux.scala 31:69:@6044.4]
  wire [15:0] _T_10354; // @[Mux.scala 31:69:@6045.4]
  wire  _T_10355; // @[OneHot.scala 66:30:@6046.4]
  wire  _T_10356; // @[OneHot.scala 66:30:@6047.4]
  wire  _T_10357; // @[OneHot.scala 66:30:@6048.4]
  wire  _T_10358; // @[OneHot.scala 66:30:@6049.4]
  wire  _T_10359; // @[OneHot.scala 66:30:@6050.4]
  wire  _T_10360; // @[OneHot.scala 66:30:@6051.4]
  wire  _T_10361; // @[OneHot.scala 66:30:@6052.4]
  wire  _T_10362; // @[OneHot.scala 66:30:@6053.4]
  wire  _T_10363; // @[OneHot.scala 66:30:@6054.4]
  wire  _T_10364; // @[OneHot.scala 66:30:@6055.4]
  wire  _T_10365; // @[OneHot.scala 66:30:@6056.4]
  wire  _T_10366; // @[OneHot.scala 66:30:@6057.4]
  wire  _T_10367; // @[OneHot.scala 66:30:@6058.4]
  wire  _T_10368; // @[OneHot.scala 66:30:@6059.4]
  wire  _T_10369; // @[OneHot.scala 66:30:@6060.4]
  wire  _T_10370; // @[OneHot.scala 66:30:@6061.4]
  wire [15:0] _T_10411; // @[Mux.scala 31:69:@6079.4]
  wire [15:0] _T_10412; // @[Mux.scala 31:69:@6080.4]
  wire [15:0] _T_10413; // @[Mux.scala 31:69:@6081.4]
  wire [15:0] _T_10414; // @[Mux.scala 31:69:@6082.4]
  wire [15:0] _T_10415; // @[Mux.scala 31:69:@6083.4]
  wire [15:0] _T_10416; // @[Mux.scala 31:69:@6084.4]
  wire [15:0] _T_10417; // @[Mux.scala 31:69:@6085.4]
  wire [15:0] _T_10418; // @[Mux.scala 31:69:@6086.4]
  wire [15:0] _T_10419; // @[Mux.scala 31:69:@6087.4]
  wire [15:0] _T_10420; // @[Mux.scala 31:69:@6088.4]
  wire [15:0] _T_10421; // @[Mux.scala 31:69:@6089.4]
  wire [15:0] _T_10422; // @[Mux.scala 31:69:@6090.4]
  wire [15:0] _T_10423; // @[Mux.scala 31:69:@6091.4]
  wire [15:0] _T_10424; // @[Mux.scala 31:69:@6092.4]
  wire [15:0] _T_10425; // @[Mux.scala 31:69:@6093.4]
  wire [15:0] _T_10426; // @[Mux.scala 31:69:@6094.4]
  wire  _T_10427; // @[OneHot.scala 66:30:@6095.4]
  wire  _T_10428; // @[OneHot.scala 66:30:@6096.4]
  wire  _T_10429; // @[OneHot.scala 66:30:@6097.4]
  wire  _T_10430; // @[OneHot.scala 66:30:@6098.4]
  wire  _T_10431; // @[OneHot.scala 66:30:@6099.4]
  wire  _T_10432; // @[OneHot.scala 66:30:@6100.4]
  wire  _T_10433; // @[OneHot.scala 66:30:@6101.4]
  wire  _T_10434; // @[OneHot.scala 66:30:@6102.4]
  wire  _T_10435; // @[OneHot.scala 66:30:@6103.4]
  wire  _T_10436; // @[OneHot.scala 66:30:@6104.4]
  wire  _T_10437; // @[OneHot.scala 66:30:@6105.4]
  wire  _T_10438; // @[OneHot.scala 66:30:@6106.4]
  wire  _T_10439; // @[OneHot.scala 66:30:@6107.4]
  wire  _T_10440; // @[OneHot.scala 66:30:@6108.4]
  wire  _T_10441; // @[OneHot.scala 66:30:@6109.4]
  wire  _T_10442; // @[OneHot.scala 66:30:@6110.4]
  wire [15:0] _T_10483; // @[Mux.scala 31:69:@6128.4]
  wire [15:0] _T_10484; // @[Mux.scala 31:69:@6129.4]
  wire [15:0] _T_10485; // @[Mux.scala 31:69:@6130.4]
  wire [15:0] _T_10486; // @[Mux.scala 31:69:@6131.4]
  wire [15:0] _T_10487; // @[Mux.scala 31:69:@6132.4]
  wire [15:0] _T_10488; // @[Mux.scala 31:69:@6133.4]
  wire [15:0] _T_10489; // @[Mux.scala 31:69:@6134.4]
  wire [15:0] _T_10490; // @[Mux.scala 31:69:@6135.4]
  wire [15:0] _T_10491; // @[Mux.scala 31:69:@6136.4]
  wire [15:0] _T_10492; // @[Mux.scala 31:69:@6137.4]
  wire [15:0] _T_10493; // @[Mux.scala 31:69:@6138.4]
  wire [15:0] _T_10494; // @[Mux.scala 31:69:@6139.4]
  wire [15:0] _T_10495; // @[Mux.scala 31:69:@6140.4]
  wire [15:0] _T_10496; // @[Mux.scala 31:69:@6141.4]
  wire [15:0] _T_10497; // @[Mux.scala 31:69:@6142.4]
  wire [15:0] _T_10498; // @[Mux.scala 31:69:@6143.4]
  wire  _T_10499; // @[OneHot.scala 66:30:@6144.4]
  wire  _T_10500; // @[OneHot.scala 66:30:@6145.4]
  wire  _T_10501; // @[OneHot.scala 66:30:@6146.4]
  wire  _T_10502; // @[OneHot.scala 66:30:@6147.4]
  wire  _T_10503; // @[OneHot.scala 66:30:@6148.4]
  wire  _T_10504; // @[OneHot.scala 66:30:@6149.4]
  wire  _T_10505; // @[OneHot.scala 66:30:@6150.4]
  wire  _T_10506; // @[OneHot.scala 66:30:@6151.4]
  wire  _T_10507; // @[OneHot.scala 66:30:@6152.4]
  wire  _T_10508; // @[OneHot.scala 66:30:@6153.4]
  wire  _T_10509; // @[OneHot.scala 66:30:@6154.4]
  wire  _T_10510; // @[OneHot.scala 66:30:@6155.4]
  wire  _T_10511; // @[OneHot.scala 66:30:@6156.4]
  wire  _T_10512; // @[OneHot.scala 66:30:@6157.4]
  wire  _T_10513; // @[OneHot.scala 66:30:@6158.4]
  wire  _T_10514; // @[OneHot.scala 66:30:@6159.4]
  wire [15:0] _T_10555; // @[Mux.scala 31:69:@6177.4]
  wire [15:0] _T_10556; // @[Mux.scala 31:69:@6178.4]
  wire [15:0] _T_10557; // @[Mux.scala 31:69:@6179.4]
  wire [15:0] _T_10558; // @[Mux.scala 31:69:@6180.4]
  wire [15:0] _T_10559; // @[Mux.scala 31:69:@6181.4]
  wire [15:0] _T_10560; // @[Mux.scala 31:69:@6182.4]
  wire [15:0] _T_10561; // @[Mux.scala 31:69:@6183.4]
  wire [15:0] _T_10562; // @[Mux.scala 31:69:@6184.4]
  wire [15:0] _T_10563; // @[Mux.scala 31:69:@6185.4]
  wire [15:0] _T_10564; // @[Mux.scala 31:69:@6186.4]
  wire [15:0] _T_10565; // @[Mux.scala 31:69:@6187.4]
  wire [15:0] _T_10566; // @[Mux.scala 31:69:@6188.4]
  wire [15:0] _T_10567; // @[Mux.scala 31:69:@6189.4]
  wire [15:0] _T_10568; // @[Mux.scala 31:69:@6190.4]
  wire [15:0] _T_10569; // @[Mux.scala 31:69:@6191.4]
  wire [15:0] _T_10570; // @[Mux.scala 31:69:@6192.4]
  wire  _T_10571; // @[OneHot.scala 66:30:@6193.4]
  wire  _T_10572; // @[OneHot.scala 66:30:@6194.4]
  wire  _T_10573; // @[OneHot.scala 66:30:@6195.4]
  wire  _T_10574; // @[OneHot.scala 66:30:@6196.4]
  wire  _T_10575; // @[OneHot.scala 66:30:@6197.4]
  wire  _T_10576; // @[OneHot.scala 66:30:@6198.4]
  wire  _T_10577; // @[OneHot.scala 66:30:@6199.4]
  wire  _T_10578; // @[OneHot.scala 66:30:@6200.4]
  wire  _T_10579; // @[OneHot.scala 66:30:@6201.4]
  wire  _T_10580; // @[OneHot.scala 66:30:@6202.4]
  wire  _T_10581; // @[OneHot.scala 66:30:@6203.4]
  wire  _T_10582; // @[OneHot.scala 66:30:@6204.4]
  wire  _T_10583; // @[OneHot.scala 66:30:@6205.4]
  wire  _T_10584; // @[OneHot.scala 66:30:@6206.4]
  wire  _T_10585; // @[OneHot.scala 66:30:@6207.4]
  wire  _T_10586; // @[OneHot.scala 66:30:@6208.4]
  wire [15:0] _T_10627; // @[Mux.scala 31:69:@6226.4]
  wire [15:0] _T_10628; // @[Mux.scala 31:69:@6227.4]
  wire [15:0] _T_10629; // @[Mux.scala 31:69:@6228.4]
  wire [15:0] _T_10630; // @[Mux.scala 31:69:@6229.4]
  wire [15:0] _T_10631; // @[Mux.scala 31:69:@6230.4]
  wire [15:0] _T_10632; // @[Mux.scala 31:69:@6231.4]
  wire [15:0] _T_10633; // @[Mux.scala 31:69:@6232.4]
  wire [15:0] _T_10634; // @[Mux.scala 31:69:@6233.4]
  wire [15:0] _T_10635; // @[Mux.scala 31:69:@6234.4]
  wire [15:0] _T_10636; // @[Mux.scala 31:69:@6235.4]
  wire [15:0] _T_10637; // @[Mux.scala 31:69:@6236.4]
  wire [15:0] _T_10638; // @[Mux.scala 31:69:@6237.4]
  wire [15:0] _T_10639; // @[Mux.scala 31:69:@6238.4]
  wire [15:0] _T_10640; // @[Mux.scala 31:69:@6239.4]
  wire [15:0] _T_10641; // @[Mux.scala 31:69:@6240.4]
  wire [15:0] _T_10642; // @[Mux.scala 31:69:@6241.4]
  wire  _T_10643; // @[OneHot.scala 66:30:@6242.4]
  wire  _T_10644; // @[OneHot.scala 66:30:@6243.4]
  wire  _T_10645; // @[OneHot.scala 66:30:@6244.4]
  wire  _T_10646; // @[OneHot.scala 66:30:@6245.4]
  wire  _T_10647; // @[OneHot.scala 66:30:@6246.4]
  wire  _T_10648; // @[OneHot.scala 66:30:@6247.4]
  wire  _T_10649; // @[OneHot.scala 66:30:@6248.4]
  wire  _T_10650; // @[OneHot.scala 66:30:@6249.4]
  wire  _T_10651; // @[OneHot.scala 66:30:@6250.4]
  wire  _T_10652; // @[OneHot.scala 66:30:@6251.4]
  wire  _T_10653; // @[OneHot.scala 66:30:@6252.4]
  wire  _T_10654; // @[OneHot.scala 66:30:@6253.4]
  wire  _T_10655; // @[OneHot.scala 66:30:@6254.4]
  wire  _T_10656; // @[OneHot.scala 66:30:@6255.4]
  wire  _T_10657; // @[OneHot.scala 66:30:@6256.4]
  wire  _T_10658; // @[OneHot.scala 66:30:@6257.4]
  wire [15:0] _T_10699; // @[Mux.scala 31:69:@6275.4]
  wire [15:0] _T_10700; // @[Mux.scala 31:69:@6276.4]
  wire [15:0] _T_10701; // @[Mux.scala 31:69:@6277.4]
  wire [15:0] _T_10702; // @[Mux.scala 31:69:@6278.4]
  wire [15:0] _T_10703; // @[Mux.scala 31:69:@6279.4]
  wire [15:0] _T_10704; // @[Mux.scala 31:69:@6280.4]
  wire [15:0] _T_10705; // @[Mux.scala 31:69:@6281.4]
  wire [15:0] _T_10706; // @[Mux.scala 31:69:@6282.4]
  wire [15:0] _T_10707; // @[Mux.scala 31:69:@6283.4]
  wire [15:0] _T_10708; // @[Mux.scala 31:69:@6284.4]
  wire [15:0] _T_10709; // @[Mux.scala 31:69:@6285.4]
  wire [15:0] _T_10710; // @[Mux.scala 31:69:@6286.4]
  wire [15:0] _T_10711; // @[Mux.scala 31:69:@6287.4]
  wire [15:0] _T_10712; // @[Mux.scala 31:69:@6288.4]
  wire [15:0] _T_10713; // @[Mux.scala 31:69:@6289.4]
  wire [15:0] _T_10714; // @[Mux.scala 31:69:@6290.4]
  wire  _T_10715; // @[OneHot.scala 66:30:@6291.4]
  wire  _T_10716; // @[OneHot.scala 66:30:@6292.4]
  wire  _T_10717; // @[OneHot.scala 66:30:@6293.4]
  wire  _T_10718; // @[OneHot.scala 66:30:@6294.4]
  wire  _T_10719; // @[OneHot.scala 66:30:@6295.4]
  wire  _T_10720; // @[OneHot.scala 66:30:@6296.4]
  wire  _T_10721; // @[OneHot.scala 66:30:@6297.4]
  wire  _T_10722; // @[OneHot.scala 66:30:@6298.4]
  wire  _T_10723; // @[OneHot.scala 66:30:@6299.4]
  wire  _T_10724; // @[OneHot.scala 66:30:@6300.4]
  wire  _T_10725; // @[OneHot.scala 66:30:@6301.4]
  wire  _T_10726; // @[OneHot.scala 66:30:@6302.4]
  wire  _T_10727; // @[OneHot.scala 66:30:@6303.4]
  wire  _T_10728; // @[OneHot.scala 66:30:@6304.4]
  wire  _T_10729; // @[OneHot.scala 66:30:@6305.4]
  wire  _T_10730; // @[OneHot.scala 66:30:@6306.4]
  wire [15:0] _T_10771; // @[Mux.scala 31:69:@6324.4]
  wire [15:0] _T_10772; // @[Mux.scala 31:69:@6325.4]
  wire [15:0] _T_10773; // @[Mux.scala 31:69:@6326.4]
  wire [15:0] _T_10774; // @[Mux.scala 31:69:@6327.4]
  wire [15:0] _T_10775; // @[Mux.scala 31:69:@6328.4]
  wire [15:0] _T_10776; // @[Mux.scala 31:69:@6329.4]
  wire [15:0] _T_10777; // @[Mux.scala 31:69:@6330.4]
  wire [15:0] _T_10778; // @[Mux.scala 31:69:@6331.4]
  wire [15:0] _T_10779; // @[Mux.scala 31:69:@6332.4]
  wire [15:0] _T_10780; // @[Mux.scala 31:69:@6333.4]
  wire [15:0] _T_10781; // @[Mux.scala 31:69:@6334.4]
  wire [15:0] _T_10782; // @[Mux.scala 31:69:@6335.4]
  wire [15:0] _T_10783; // @[Mux.scala 31:69:@6336.4]
  wire [15:0] _T_10784; // @[Mux.scala 31:69:@6337.4]
  wire [15:0] _T_10785; // @[Mux.scala 31:69:@6338.4]
  wire [15:0] _T_10786; // @[Mux.scala 31:69:@6339.4]
  wire  _T_10787; // @[OneHot.scala 66:30:@6340.4]
  wire  _T_10788; // @[OneHot.scala 66:30:@6341.4]
  wire  _T_10789; // @[OneHot.scala 66:30:@6342.4]
  wire  _T_10790; // @[OneHot.scala 66:30:@6343.4]
  wire  _T_10791; // @[OneHot.scala 66:30:@6344.4]
  wire  _T_10792; // @[OneHot.scala 66:30:@6345.4]
  wire  _T_10793; // @[OneHot.scala 66:30:@6346.4]
  wire  _T_10794; // @[OneHot.scala 66:30:@6347.4]
  wire  _T_10795; // @[OneHot.scala 66:30:@6348.4]
  wire  _T_10796; // @[OneHot.scala 66:30:@6349.4]
  wire  _T_10797; // @[OneHot.scala 66:30:@6350.4]
  wire  _T_10798; // @[OneHot.scala 66:30:@6351.4]
  wire  _T_10799; // @[OneHot.scala 66:30:@6352.4]
  wire  _T_10800; // @[OneHot.scala 66:30:@6353.4]
  wire  _T_10801; // @[OneHot.scala 66:30:@6354.4]
  wire  _T_10802; // @[OneHot.scala 66:30:@6355.4]
  wire [7:0] _T_10867; // @[Mux.scala 19:72:@6379.4]
  wire [15:0] _T_10875; // @[Mux.scala 19:72:@6387.4]
  wire [15:0] _T_10877; // @[Mux.scala 19:72:@6388.4]
  wire [7:0] _T_10884; // @[Mux.scala 19:72:@6395.4]
  wire [15:0] _T_10892; // @[Mux.scala 19:72:@6403.4]
  wire [15:0] _T_10894; // @[Mux.scala 19:72:@6404.4]
  wire [7:0] _T_10901; // @[Mux.scala 19:72:@6411.4]
  wire [15:0] _T_10909; // @[Mux.scala 19:72:@6419.4]
  wire [15:0] _T_10911; // @[Mux.scala 19:72:@6420.4]
  wire [7:0] _T_10918; // @[Mux.scala 19:72:@6427.4]
  wire [15:0] _T_10926; // @[Mux.scala 19:72:@6435.4]
  wire [15:0] _T_10928; // @[Mux.scala 19:72:@6436.4]
  wire [7:0] _T_10935; // @[Mux.scala 19:72:@6443.4]
  wire [15:0] _T_10943; // @[Mux.scala 19:72:@6451.4]
  wire [15:0] _T_10945; // @[Mux.scala 19:72:@6452.4]
  wire [7:0] _T_10952; // @[Mux.scala 19:72:@6459.4]
  wire [15:0] _T_10960; // @[Mux.scala 19:72:@6467.4]
  wire [15:0] _T_10962; // @[Mux.scala 19:72:@6468.4]
  wire [7:0] _T_10969; // @[Mux.scala 19:72:@6475.4]
  wire [15:0] _T_10977; // @[Mux.scala 19:72:@6483.4]
  wire [15:0] _T_10979; // @[Mux.scala 19:72:@6484.4]
  wire [7:0] _T_10986; // @[Mux.scala 19:72:@6491.4]
  wire [15:0] _T_10994; // @[Mux.scala 19:72:@6499.4]
  wire [15:0] _T_10996; // @[Mux.scala 19:72:@6500.4]
  wire [7:0] _T_11003; // @[Mux.scala 19:72:@6507.4]
  wire [15:0] _T_11011; // @[Mux.scala 19:72:@6515.4]
  wire [15:0] _T_11013; // @[Mux.scala 19:72:@6516.4]
  wire [7:0] _T_11020; // @[Mux.scala 19:72:@6523.4]
  wire [15:0] _T_11028; // @[Mux.scala 19:72:@6531.4]
  wire [15:0] _T_11030; // @[Mux.scala 19:72:@6532.4]
  wire [7:0] _T_11037; // @[Mux.scala 19:72:@6539.4]
  wire [15:0] _T_11045; // @[Mux.scala 19:72:@6547.4]
  wire [15:0] _T_11047; // @[Mux.scala 19:72:@6548.4]
  wire [7:0] _T_11054; // @[Mux.scala 19:72:@6555.4]
  wire [15:0] _T_11062; // @[Mux.scala 19:72:@6563.4]
  wire [15:0] _T_11064; // @[Mux.scala 19:72:@6564.4]
  wire [7:0] _T_11071; // @[Mux.scala 19:72:@6571.4]
  wire [15:0] _T_11079; // @[Mux.scala 19:72:@6579.4]
  wire [15:0] _T_11081; // @[Mux.scala 19:72:@6580.4]
  wire [7:0] _T_11088; // @[Mux.scala 19:72:@6587.4]
  wire [15:0] _T_11096; // @[Mux.scala 19:72:@6595.4]
  wire [15:0] _T_11098; // @[Mux.scala 19:72:@6596.4]
  wire [7:0] _T_11105; // @[Mux.scala 19:72:@6603.4]
  wire [15:0] _T_11113; // @[Mux.scala 19:72:@6611.4]
  wire [15:0] _T_11115; // @[Mux.scala 19:72:@6612.4]
  wire [7:0] _T_11122; // @[Mux.scala 19:72:@6619.4]
  wire [15:0] _T_11130; // @[Mux.scala 19:72:@6627.4]
  wire [15:0] _T_11132; // @[Mux.scala 19:72:@6628.4]
  wire [15:0] _T_11133; // @[Mux.scala 19:72:@6629.4]
  wire [15:0] _T_11134; // @[Mux.scala 19:72:@6630.4]
  wire [15:0] _T_11135; // @[Mux.scala 19:72:@6631.4]
  wire [15:0] _T_11136; // @[Mux.scala 19:72:@6632.4]
  wire [15:0] _T_11137; // @[Mux.scala 19:72:@6633.4]
  wire [15:0] _T_11138; // @[Mux.scala 19:72:@6634.4]
  wire [15:0] _T_11139; // @[Mux.scala 19:72:@6635.4]
  wire [15:0] _T_11140; // @[Mux.scala 19:72:@6636.4]
  wire [15:0] _T_11141; // @[Mux.scala 19:72:@6637.4]
  wire [15:0] _T_11142; // @[Mux.scala 19:72:@6638.4]
  wire [15:0] _T_11143; // @[Mux.scala 19:72:@6639.4]
  wire [15:0] _T_11144; // @[Mux.scala 19:72:@6640.4]
  wire [15:0] _T_11145; // @[Mux.scala 19:72:@6641.4]
  wire [15:0] _T_11146; // @[Mux.scala 19:72:@6642.4]
  wire [15:0] _T_11147; // @[Mux.scala 19:72:@6643.4]
  wire  inputDataPriorityPorts_1_0; // @[Mux.scala 19:72:@6647.4]
  wire  inputDataPriorityPorts_1_1; // @[Mux.scala 19:72:@6649.4]
  wire  inputDataPriorityPorts_1_2; // @[Mux.scala 19:72:@6651.4]
  wire  inputDataPriorityPorts_1_3; // @[Mux.scala 19:72:@6653.4]
  wire  inputDataPriorityPorts_1_4; // @[Mux.scala 19:72:@6655.4]
  wire  inputDataPriorityPorts_1_5; // @[Mux.scala 19:72:@6657.4]
  wire  inputDataPriorityPorts_1_6; // @[Mux.scala 19:72:@6659.4]
  wire  inputDataPriorityPorts_1_7; // @[Mux.scala 19:72:@6661.4]
  wire  inputDataPriorityPorts_1_8; // @[Mux.scala 19:72:@6663.4]
  wire  inputDataPriorityPorts_1_9; // @[Mux.scala 19:72:@6665.4]
  wire  inputDataPriorityPorts_1_10; // @[Mux.scala 19:72:@6667.4]
  wire  inputDataPriorityPorts_1_11; // @[Mux.scala 19:72:@6669.4]
  wire  inputDataPriorityPorts_1_12; // @[Mux.scala 19:72:@6671.4]
  wire  inputDataPriorityPorts_1_13; // @[Mux.scala 19:72:@6673.4]
  wire  inputDataPriorityPorts_1_14; // @[Mux.scala 19:72:@6675.4]
  wire  inputDataPriorityPorts_1_15; // @[Mux.scala 19:72:@6677.4]
  wire  _T_11293; // @[StoreQueue.scala 209:52:@6701.6]
  wire  _T_11294; // @[StoreQueue.scala 209:81:@6702.6]
  wire  _T_11297; // @[StoreQueue.scala 209:52:@6704.6]
  wire  _T_11298; // @[StoreQueue.scala 209:81:@6705.6]
  wire  _T_11309; // @[StoreQueue.scala 210:30:@6710.6]
  wire [1:0] _T_11310; // @[OneHot.scala 18:45:@6712.8]
  wire  _T_11311; // @[CircuitMath.scala 30:8:@6713.8]
  wire [31:0] _GEN_993; // @[StoreQueue.scala 211:30:@6714.8]
  wire [31:0] _GEN_994; // @[StoreQueue.scala 210:40:@6711.6]
  wire  _GEN_995; // @[StoreQueue.scala 210:40:@6711.6]
  wire  _T_11316; // @[StoreQueue.scala 215:52:@6718.6]
  wire  _T_11317; // @[StoreQueue.scala 215:81:@6719.6]
  wire  _T_11320; // @[StoreQueue.scala 215:52:@6721.6]
  wire  _T_11321; // @[StoreQueue.scala 215:81:@6722.6]
  wire  _T_11332; // @[StoreQueue.scala 216:30:@6727.6]
  wire [1:0] _T_11333; // @[OneHot.scala 18:45:@6729.8]
  wire  _T_11334; // @[CircuitMath.scala 30:8:@6730.8]
  wire [31:0] _GEN_997; // @[StoreQueue.scala 217:30:@6731.8]
  wire [31:0] _GEN_998; // @[StoreQueue.scala 216:40:@6728.6]
  wire  _GEN_999; // @[StoreQueue.scala 216:40:@6728.6]
  wire  _GEN_1000; // @[StoreQueue.scala 204:35:@6695.4]
  wire  _GEN_1001; // @[StoreQueue.scala 204:35:@6695.4]
  wire [31:0] _GEN_1002; // @[StoreQueue.scala 204:35:@6695.4]
  wire [31:0] _GEN_1003; // @[StoreQueue.scala 204:35:@6695.4]
  wire  _T_11341; // @[StoreQueue.scala 209:52:@6741.6]
  wire  _T_11342; // @[StoreQueue.scala 209:81:@6742.6]
  wire  _T_11345; // @[StoreQueue.scala 209:52:@6744.6]
  wire  _T_11346; // @[StoreQueue.scala 209:81:@6745.6]
  wire  _T_11357; // @[StoreQueue.scala 210:30:@6750.6]
  wire [1:0] _T_11358; // @[OneHot.scala 18:45:@6752.8]
  wire  _T_11359; // @[CircuitMath.scala 30:8:@6753.8]
  wire [31:0] _GEN_1005; // @[StoreQueue.scala 211:30:@6754.8]
  wire [31:0] _GEN_1006; // @[StoreQueue.scala 210:40:@6751.6]
  wire  _GEN_1007; // @[StoreQueue.scala 210:40:@6751.6]
  wire  _T_11364; // @[StoreQueue.scala 215:52:@6758.6]
  wire  _T_11365; // @[StoreQueue.scala 215:81:@6759.6]
  wire  _T_11368; // @[StoreQueue.scala 215:52:@6761.6]
  wire  _T_11369; // @[StoreQueue.scala 215:81:@6762.6]
  wire  _T_11380; // @[StoreQueue.scala 216:30:@6767.6]
  wire [1:0] _T_11381; // @[OneHot.scala 18:45:@6769.8]
  wire  _T_11382; // @[CircuitMath.scala 30:8:@6770.8]
  wire [31:0] _GEN_1009; // @[StoreQueue.scala 217:30:@6771.8]
  wire [31:0] _GEN_1010; // @[StoreQueue.scala 216:40:@6768.6]
  wire  _GEN_1011; // @[StoreQueue.scala 216:40:@6768.6]
  wire  _GEN_1012; // @[StoreQueue.scala 204:35:@6735.4]
  wire  _GEN_1013; // @[StoreQueue.scala 204:35:@6735.4]
  wire [31:0] _GEN_1014; // @[StoreQueue.scala 204:35:@6735.4]
  wire [31:0] _GEN_1015; // @[StoreQueue.scala 204:35:@6735.4]
  wire  _T_11389; // @[StoreQueue.scala 209:52:@6781.6]
  wire  _T_11390; // @[StoreQueue.scala 209:81:@6782.6]
  wire  _T_11393; // @[StoreQueue.scala 209:52:@6784.6]
  wire  _T_11394; // @[StoreQueue.scala 209:81:@6785.6]
  wire  _T_11405; // @[StoreQueue.scala 210:30:@6790.6]
  wire [1:0] _T_11406; // @[OneHot.scala 18:45:@6792.8]
  wire  _T_11407; // @[CircuitMath.scala 30:8:@6793.8]
  wire [31:0] _GEN_1017; // @[StoreQueue.scala 211:30:@6794.8]
  wire [31:0] _GEN_1018; // @[StoreQueue.scala 210:40:@6791.6]
  wire  _GEN_1019; // @[StoreQueue.scala 210:40:@6791.6]
  wire  _T_11412; // @[StoreQueue.scala 215:52:@6798.6]
  wire  _T_11413; // @[StoreQueue.scala 215:81:@6799.6]
  wire  _T_11416; // @[StoreQueue.scala 215:52:@6801.6]
  wire  _T_11417; // @[StoreQueue.scala 215:81:@6802.6]
  wire  _T_11428; // @[StoreQueue.scala 216:30:@6807.6]
  wire [1:0] _T_11429; // @[OneHot.scala 18:45:@6809.8]
  wire  _T_11430; // @[CircuitMath.scala 30:8:@6810.8]
  wire [31:0] _GEN_1021; // @[StoreQueue.scala 217:30:@6811.8]
  wire [31:0] _GEN_1022; // @[StoreQueue.scala 216:40:@6808.6]
  wire  _GEN_1023; // @[StoreQueue.scala 216:40:@6808.6]
  wire  _GEN_1024; // @[StoreQueue.scala 204:35:@6775.4]
  wire  _GEN_1025; // @[StoreQueue.scala 204:35:@6775.4]
  wire [31:0] _GEN_1026; // @[StoreQueue.scala 204:35:@6775.4]
  wire [31:0] _GEN_1027; // @[StoreQueue.scala 204:35:@6775.4]
  wire  _T_11437; // @[StoreQueue.scala 209:52:@6821.6]
  wire  _T_11438; // @[StoreQueue.scala 209:81:@6822.6]
  wire  _T_11441; // @[StoreQueue.scala 209:52:@6824.6]
  wire  _T_11442; // @[StoreQueue.scala 209:81:@6825.6]
  wire  _T_11453; // @[StoreQueue.scala 210:30:@6830.6]
  wire [1:0] _T_11454; // @[OneHot.scala 18:45:@6832.8]
  wire  _T_11455; // @[CircuitMath.scala 30:8:@6833.8]
  wire [31:0] _GEN_1029; // @[StoreQueue.scala 211:30:@6834.8]
  wire [31:0] _GEN_1030; // @[StoreQueue.scala 210:40:@6831.6]
  wire  _GEN_1031; // @[StoreQueue.scala 210:40:@6831.6]
  wire  _T_11460; // @[StoreQueue.scala 215:52:@6838.6]
  wire  _T_11461; // @[StoreQueue.scala 215:81:@6839.6]
  wire  _T_11464; // @[StoreQueue.scala 215:52:@6841.6]
  wire  _T_11465; // @[StoreQueue.scala 215:81:@6842.6]
  wire  _T_11476; // @[StoreQueue.scala 216:30:@6847.6]
  wire [1:0] _T_11477; // @[OneHot.scala 18:45:@6849.8]
  wire  _T_11478; // @[CircuitMath.scala 30:8:@6850.8]
  wire [31:0] _GEN_1033; // @[StoreQueue.scala 217:30:@6851.8]
  wire [31:0] _GEN_1034; // @[StoreQueue.scala 216:40:@6848.6]
  wire  _GEN_1035; // @[StoreQueue.scala 216:40:@6848.6]
  wire  _GEN_1036; // @[StoreQueue.scala 204:35:@6815.4]
  wire  _GEN_1037; // @[StoreQueue.scala 204:35:@6815.4]
  wire [31:0] _GEN_1038; // @[StoreQueue.scala 204:35:@6815.4]
  wire [31:0] _GEN_1039; // @[StoreQueue.scala 204:35:@6815.4]
  wire  _T_11485; // @[StoreQueue.scala 209:52:@6861.6]
  wire  _T_11486; // @[StoreQueue.scala 209:81:@6862.6]
  wire  _T_11489; // @[StoreQueue.scala 209:52:@6864.6]
  wire  _T_11490; // @[StoreQueue.scala 209:81:@6865.6]
  wire  _T_11501; // @[StoreQueue.scala 210:30:@6870.6]
  wire [1:0] _T_11502; // @[OneHot.scala 18:45:@6872.8]
  wire  _T_11503; // @[CircuitMath.scala 30:8:@6873.8]
  wire [31:0] _GEN_1041; // @[StoreQueue.scala 211:30:@6874.8]
  wire [31:0] _GEN_1042; // @[StoreQueue.scala 210:40:@6871.6]
  wire  _GEN_1043; // @[StoreQueue.scala 210:40:@6871.6]
  wire  _T_11508; // @[StoreQueue.scala 215:52:@6878.6]
  wire  _T_11509; // @[StoreQueue.scala 215:81:@6879.6]
  wire  _T_11512; // @[StoreQueue.scala 215:52:@6881.6]
  wire  _T_11513; // @[StoreQueue.scala 215:81:@6882.6]
  wire  _T_11524; // @[StoreQueue.scala 216:30:@6887.6]
  wire [1:0] _T_11525; // @[OneHot.scala 18:45:@6889.8]
  wire  _T_11526; // @[CircuitMath.scala 30:8:@6890.8]
  wire [31:0] _GEN_1045; // @[StoreQueue.scala 217:30:@6891.8]
  wire [31:0] _GEN_1046; // @[StoreQueue.scala 216:40:@6888.6]
  wire  _GEN_1047; // @[StoreQueue.scala 216:40:@6888.6]
  wire  _GEN_1048; // @[StoreQueue.scala 204:35:@6855.4]
  wire  _GEN_1049; // @[StoreQueue.scala 204:35:@6855.4]
  wire [31:0] _GEN_1050; // @[StoreQueue.scala 204:35:@6855.4]
  wire [31:0] _GEN_1051; // @[StoreQueue.scala 204:35:@6855.4]
  wire  _T_11533; // @[StoreQueue.scala 209:52:@6901.6]
  wire  _T_11534; // @[StoreQueue.scala 209:81:@6902.6]
  wire  _T_11537; // @[StoreQueue.scala 209:52:@6904.6]
  wire  _T_11538; // @[StoreQueue.scala 209:81:@6905.6]
  wire  _T_11549; // @[StoreQueue.scala 210:30:@6910.6]
  wire [1:0] _T_11550; // @[OneHot.scala 18:45:@6912.8]
  wire  _T_11551; // @[CircuitMath.scala 30:8:@6913.8]
  wire [31:0] _GEN_1053; // @[StoreQueue.scala 211:30:@6914.8]
  wire [31:0] _GEN_1054; // @[StoreQueue.scala 210:40:@6911.6]
  wire  _GEN_1055; // @[StoreQueue.scala 210:40:@6911.6]
  wire  _T_11556; // @[StoreQueue.scala 215:52:@6918.6]
  wire  _T_11557; // @[StoreQueue.scala 215:81:@6919.6]
  wire  _T_11560; // @[StoreQueue.scala 215:52:@6921.6]
  wire  _T_11561; // @[StoreQueue.scala 215:81:@6922.6]
  wire  _T_11572; // @[StoreQueue.scala 216:30:@6927.6]
  wire [1:0] _T_11573; // @[OneHot.scala 18:45:@6929.8]
  wire  _T_11574; // @[CircuitMath.scala 30:8:@6930.8]
  wire [31:0] _GEN_1057; // @[StoreQueue.scala 217:30:@6931.8]
  wire [31:0] _GEN_1058; // @[StoreQueue.scala 216:40:@6928.6]
  wire  _GEN_1059; // @[StoreQueue.scala 216:40:@6928.6]
  wire  _GEN_1060; // @[StoreQueue.scala 204:35:@6895.4]
  wire  _GEN_1061; // @[StoreQueue.scala 204:35:@6895.4]
  wire [31:0] _GEN_1062; // @[StoreQueue.scala 204:35:@6895.4]
  wire [31:0] _GEN_1063; // @[StoreQueue.scala 204:35:@6895.4]
  wire  _T_11581; // @[StoreQueue.scala 209:52:@6941.6]
  wire  _T_11582; // @[StoreQueue.scala 209:81:@6942.6]
  wire  _T_11585; // @[StoreQueue.scala 209:52:@6944.6]
  wire  _T_11586; // @[StoreQueue.scala 209:81:@6945.6]
  wire  _T_11597; // @[StoreQueue.scala 210:30:@6950.6]
  wire [1:0] _T_11598; // @[OneHot.scala 18:45:@6952.8]
  wire  _T_11599; // @[CircuitMath.scala 30:8:@6953.8]
  wire [31:0] _GEN_1065; // @[StoreQueue.scala 211:30:@6954.8]
  wire [31:0] _GEN_1066; // @[StoreQueue.scala 210:40:@6951.6]
  wire  _GEN_1067; // @[StoreQueue.scala 210:40:@6951.6]
  wire  _T_11604; // @[StoreQueue.scala 215:52:@6958.6]
  wire  _T_11605; // @[StoreQueue.scala 215:81:@6959.6]
  wire  _T_11608; // @[StoreQueue.scala 215:52:@6961.6]
  wire  _T_11609; // @[StoreQueue.scala 215:81:@6962.6]
  wire  _T_11620; // @[StoreQueue.scala 216:30:@6967.6]
  wire [1:0] _T_11621; // @[OneHot.scala 18:45:@6969.8]
  wire  _T_11622; // @[CircuitMath.scala 30:8:@6970.8]
  wire [31:0] _GEN_1069; // @[StoreQueue.scala 217:30:@6971.8]
  wire [31:0] _GEN_1070; // @[StoreQueue.scala 216:40:@6968.6]
  wire  _GEN_1071; // @[StoreQueue.scala 216:40:@6968.6]
  wire  _GEN_1072; // @[StoreQueue.scala 204:35:@6935.4]
  wire  _GEN_1073; // @[StoreQueue.scala 204:35:@6935.4]
  wire [31:0] _GEN_1074; // @[StoreQueue.scala 204:35:@6935.4]
  wire [31:0] _GEN_1075; // @[StoreQueue.scala 204:35:@6935.4]
  wire  _T_11629; // @[StoreQueue.scala 209:52:@6981.6]
  wire  _T_11630; // @[StoreQueue.scala 209:81:@6982.6]
  wire  _T_11633; // @[StoreQueue.scala 209:52:@6984.6]
  wire  _T_11634; // @[StoreQueue.scala 209:81:@6985.6]
  wire  _T_11645; // @[StoreQueue.scala 210:30:@6990.6]
  wire [1:0] _T_11646; // @[OneHot.scala 18:45:@6992.8]
  wire  _T_11647; // @[CircuitMath.scala 30:8:@6993.8]
  wire [31:0] _GEN_1077; // @[StoreQueue.scala 211:30:@6994.8]
  wire [31:0] _GEN_1078; // @[StoreQueue.scala 210:40:@6991.6]
  wire  _GEN_1079; // @[StoreQueue.scala 210:40:@6991.6]
  wire  _T_11652; // @[StoreQueue.scala 215:52:@6998.6]
  wire  _T_11653; // @[StoreQueue.scala 215:81:@6999.6]
  wire  _T_11656; // @[StoreQueue.scala 215:52:@7001.6]
  wire  _T_11657; // @[StoreQueue.scala 215:81:@7002.6]
  wire  _T_11668; // @[StoreQueue.scala 216:30:@7007.6]
  wire [1:0] _T_11669; // @[OneHot.scala 18:45:@7009.8]
  wire  _T_11670; // @[CircuitMath.scala 30:8:@7010.8]
  wire [31:0] _GEN_1081; // @[StoreQueue.scala 217:30:@7011.8]
  wire [31:0] _GEN_1082; // @[StoreQueue.scala 216:40:@7008.6]
  wire  _GEN_1083; // @[StoreQueue.scala 216:40:@7008.6]
  wire  _GEN_1084; // @[StoreQueue.scala 204:35:@6975.4]
  wire  _GEN_1085; // @[StoreQueue.scala 204:35:@6975.4]
  wire [31:0] _GEN_1086; // @[StoreQueue.scala 204:35:@6975.4]
  wire [31:0] _GEN_1087; // @[StoreQueue.scala 204:35:@6975.4]
  wire  _T_11677; // @[StoreQueue.scala 209:52:@7021.6]
  wire  _T_11678; // @[StoreQueue.scala 209:81:@7022.6]
  wire  _T_11681; // @[StoreQueue.scala 209:52:@7024.6]
  wire  _T_11682; // @[StoreQueue.scala 209:81:@7025.6]
  wire  _T_11693; // @[StoreQueue.scala 210:30:@7030.6]
  wire [1:0] _T_11694; // @[OneHot.scala 18:45:@7032.8]
  wire  _T_11695; // @[CircuitMath.scala 30:8:@7033.8]
  wire [31:0] _GEN_1089; // @[StoreQueue.scala 211:30:@7034.8]
  wire [31:0] _GEN_1090; // @[StoreQueue.scala 210:40:@7031.6]
  wire  _GEN_1091; // @[StoreQueue.scala 210:40:@7031.6]
  wire  _T_11700; // @[StoreQueue.scala 215:52:@7038.6]
  wire  _T_11701; // @[StoreQueue.scala 215:81:@7039.6]
  wire  _T_11704; // @[StoreQueue.scala 215:52:@7041.6]
  wire  _T_11705; // @[StoreQueue.scala 215:81:@7042.6]
  wire  _T_11716; // @[StoreQueue.scala 216:30:@7047.6]
  wire [1:0] _T_11717; // @[OneHot.scala 18:45:@7049.8]
  wire  _T_11718; // @[CircuitMath.scala 30:8:@7050.8]
  wire [31:0] _GEN_1093; // @[StoreQueue.scala 217:30:@7051.8]
  wire [31:0] _GEN_1094; // @[StoreQueue.scala 216:40:@7048.6]
  wire  _GEN_1095; // @[StoreQueue.scala 216:40:@7048.6]
  wire  _GEN_1096; // @[StoreQueue.scala 204:35:@7015.4]
  wire  _GEN_1097; // @[StoreQueue.scala 204:35:@7015.4]
  wire [31:0] _GEN_1098; // @[StoreQueue.scala 204:35:@7015.4]
  wire [31:0] _GEN_1099; // @[StoreQueue.scala 204:35:@7015.4]
  wire  _T_11725; // @[StoreQueue.scala 209:52:@7061.6]
  wire  _T_11726; // @[StoreQueue.scala 209:81:@7062.6]
  wire  _T_11729; // @[StoreQueue.scala 209:52:@7064.6]
  wire  _T_11730; // @[StoreQueue.scala 209:81:@7065.6]
  wire  _T_11741; // @[StoreQueue.scala 210:30:@7070.6]
  wire [1:0] _T_11742; // @[OneHot.scala 18:45:@7072.8]
  wire  _T_11743; // @[CircuitMath.scala 30:8:@7073.8]
  wire [31:0] _GEN_1101; // @[StoreQueue.scala 211:30:@7074.8]
  wire [31:0] _GEN_1102; // @[StoreQueue.scala 210:40:@7071.6]
  wire  _GEN_1103; // @[StoreQueue.scala 210:40:@7071.6]
  wire  _T_11748; // @[StoreQueue.scala 215:52:@7078.6]
  wire  _T_11749; // @[StoreQueue.scala 215:81:@7079.6]
  wire  _T_11752; // @[StoreQueue.scala 215:52:@7081.6]
  wire  _T_11753; // @[StoreQueue.scala 215:81:@7082.6]
  wire  _T_11764; // @[StoreQueue.scala 216:30:@7087.6]
  wire [1:0] _T_11765; // @[OneHot.scala 18:45:@7089.8]
  wire  _T_11766; // @[CircuitMath.scala 30:8:@7090.8]
  wire [31:0] _GEN_1105; // @[StoreQueue.scala 217:30:@7091.8]
  wire [31:0] _GEN_1106; // @[StoreQueue.scala 216:40:@7088.6]
  wire  _GEN_1107; // @[StoreQueue.scala 216:40:@7088.6]
  wire  _GEN_1108; // @[StoreQueue.scala 204:35:@7055.4]
  wire  _GEN_1109; // @[StoreQueue.scala 204:35:@7055.4]
  wire [31:0] _GEN_1110; // @[StoreQueue.scala 204:35:@7055.4]
  wire [31:0] _GEN_1111; // @[StoreQueue.scala 204:35:@7055.4]
  wire  _T_11773; // @[StoreQueue.scala 209:52:@7101.6]
  wire  _T_11774; // @[StoreQueue.scala 209:81:@7102.6]
  wire  _T_11777; // @[StoreQueue.scala 209:52:@7104.6]
  wire  _T_11778; // @[StoreQueue.scala 209:81:@7105.6]
  wire  _T_11789; // @[StoreQueue.scala 210:30:@7110.6]
  wire [1:0] _T_11790; // @[OneHot.scala 18:45:@7112.8]
  wire  _T_11791; // @[CircuitMath.scala 30:8:@7113.8]
  wire [31:0] _GEN_1113; // @[StoreQueue.scala 211:30:@7114.8]
  wire [31:0] _GEN_1114; // @[StoreQueue.scala 210:40:@7111.6]
  wire  _GEN_1115; // @[StoreQueue.scala 210:40:@7111.6]
  wire  _T_11796; // @[StoreQueue.scala 215:52:@7118.6]
  wire  _T_11797; // @[StoreQueue.scala 215:81:@7119.6]
  wire  _T_11800; // @[StoreQueue.scala 215:52:@7121.6]
  wire  _T_11801; // @[StoreQueue.scala 215:81:@7122.6]
  wire  _T_11812; // @[StoreQueue.scala 216:30:@7127.6]
  wire [1:0] _T_11813; // @[OneHot.scala 18:45:@7129.8]
  wire  _T_11814; // @[CircuitMath.scala 30:8:@7130.8]
  wire [31:0] _GEN_1117; // @[StoreQueue.scala 217:30:@7131.8]
  wire [31:0] _GEN_1118; // @[StoreQueue.scala 216:40:@7128.6]
  wire  _GEN_1119; // @[StoreQueue.scala 216:40:@7128.6]
  wire  _GEN_1120; // @[StoreQueue.scala 204:35:@7095.4]
  wire  _GEN_1121; // @[StoreQueue.scala 204:35:@7095.4]
  wire [31:0] _GEN_1122; // @[StoreQueue.scala 204:35:@7095.4]
  wire [31:0] _GEN_1123; // @[StoreQueue.scala 204:35:@7095.4]
  wire  _T_11821; // @[StoreQueue.scala 209:52:@7141.6]
  wire  _T_11822; // @[StoreQueue.scala 209:81:@7142.6]
  wire  _T_11825; // @[StoreQueue.scala 209:52:@7144.6]
  wire  _T_11826; // @[StoreQueue.scala 209:81:@7145.6]
  wire  _T_11837; // @[StoreQueue.scala 210:30:@7150.6]
  wire [1:0] _T_11838; // @[OneHot.scala 18:45:@7152.8]
  wire  _T_11839; // @[CircuitMath.scala 30:8:@7153.8]
  wire [31:0] _GEN_1125; // @[StoreQueue.scala 211:30:@7154.8]
  wire [31:0] _GEN_1126; // @[StoreQueue.scala 210:40:@7151.6]
  wire  _GEN_1127; // @[StoreQueue.scala 210:40:@7151.6]
  wire  _T_11844; // @[StoreQueue.scala 215:52:@7158.6]
  wire  _T_11845; // @[StoreQueue.scala 215:81:@7159.6]
  wire  _T_11848; // @[StoreQueue.scala 215:52:@7161.6]
  wire  _T_11849; // @[StoreQueue.scala 215:81:@7162.6]
  wire  _T_11860; // @[StoreQueue.scala 216:30:@7167.6]
  wire [1:0] _T_11861; // @[OneHot.scala 18:45:@7169.8]
  wire  _T_11862; // @[CircuitMath.scala 30:8:@7170.8]
  wire [31:0] _GEN_1129; // @[StoreQueue.scala 217:30:@7171.8]
  wire [31:0] _GEN_1130; // @[StoreQueue.scala 216:40:@7168.6]
  wire  _GEN_1131; // @[StoreQueue.scala 216:40:@7168.6]
  wire  _GEN_1132; // @[StoreQueue.scala 204:35:@7135.4]
  wire  _GEN_1133; // @[StoreQueue.scala 204:35:@7135.4]
  wire [31:0] _GEN_1134; // @[StoreQueue.scala 204:35:@7135.4]
  wire [31:0] _GEN_1135; // @[StoreQueue.scala 204:35:@7135.4]
  wire  _T_11869; // @[StoreQueue.scala 209:52:@7181.6]
  wire  _T_11870; // @[StoreQueue.scala 209:81:@7182.6]
  wire  _T_11873; // @[StoreQueue.scala 209:52:@7184.6]
  wire  _T_11874; // @[StoreQueue.scala 209:81:@7185.6]
  wire  _T_11885; // @[StoreQueue.scala 210:30:@7190.6]
  wire [1:0] _T_11886; // @[OneHot.scala 18:45:@7192.8]
  wire  _T_11887; // @[CircuitMath.scala 30:8:@7193.8]
  wire [31:0] _GEN_1137; // @[StoreQueue.scala 211:30:@7194.8]
  wire [31:0] _GEN_1138; // @[StoreQueue.scala 210:40:@7191.6]
  wire  _GEN_1139; // @[StoreQueue.scala 210:40:@7191.6]
  wire  _T_11892; // @[StoreQueue.scala 215:52:@7198.6]
  wire  _T_11893; // @[StoreQueue.scala 215:81:@7199.6]
  wire  _T_11896; // @[StoreQueue.scala 215:52:@7201.6]
  wire  _T_11897; // @[StoreQueue.scala 215:81:@7202.6]
  wire  _T_11908; // @[StoreQueue.scala 216:30:@7207.6]
  wire [1:0] _T_11909; // @[OneHot.scala 18:45:@7209.8]
  wire  _T_11910; // @[CircuitMath.scala 30:8:@7210.8]
  wire [31:0] _GEN_1141; // @[StoreQueue.scala 217:30:@7211.8]
  wire [31:0] _GEN_1142; // @[StoreQueue.scala 216:40:@7208.6]
  wire  _GEN_1143; // @[StoreQueue.scala 216:40:@7208.6]
  wire  _GEN_1144; // @[StoreQueue.scala 204:35:@7175.4]
  wire  _GEN_1145; // @[StoreQueue.scala 204:35:@7175.4]
  wire [31:0] _GEN_1146; // @[StoreQueue.scala 204:35:@7175.4]
  wire [31:0] _GEN_1147; // @[StoreQueue.scala 204:35:@7175.4]
  wire  _T_11917; // @[StoreQueue.scala 209:52:@7221.6]
  wire  _T_11918; // @[StoreQueue.scala 209:81:@7222.6]
  wire  _T_11921; // @[StoreQueue.scala 209:52:@7224.6]
  wire  _T_11922; // @[StoreQueue.scala 209:81:@7225.6]
  wire  _T_11933; // @[StoreQueue.scala 210:30:@7230.6]
  wire [1:0] _T_11934; // @[OneHot.scala 18:45:@7232.8]
  wire  _T_11935; // @[CircuitMath.scala 30:8:@7233.8]
  wire [31:0] _GEN_1149; // @[StoreQueue.scala 211:30:@7234.8]
  wire [31:0] _GEN_1150; // @[StoreQueue.scala 210:40:@7231.6]
  wire  _GEN_1151; // @[StoreQueue.scala 210:40:@7231.6]
  wire  _T_11940; // @[StoreQueue.scala 215:52:@7238.6]
  wire  _T_11941; // @[StoreQueue.scala 215:81:@7239.6]
  wire  _T_11944; // @[StoreQueue.scala 215:52:@7241.6]
  wire  _T_11945; // @[StoreQueue.scala 215:81:@7242.6]
  wire  _T_11956; // @[StoreQueue.scala 216:30:@7247.6]
  wire [1:0] _T_11957; // @[OneHot.scala 18:45:@7249.8]
  wire  _T_11958; // @[CircuitMath.scala 30:8:@7250.8]
  wire [31:0] _GEN_1153; // @[StoreQueue.scala 217:30:@7251.8]
  wire [31:0] _GEN_1154; // @[StoreQueue.scala 216:40:@7248.6]
  wire  _GEN_1155; // @[StoreQueue.scala 216:40:@7248.6]
  wire  _GEN_1156; // @[StoreQueue.scala 204:35:@7215.4]
  wire  _GEN_1157; // @[StoreQueue.scala 204:35:@7215.4]
  wire [31:0] _GEN_1158; // @[StoreQueue.scala 204:35:@7215.4]
  wire [31:0] _GEN_1159; // @[StoreQueue.scala 204:35:@7215.4]
  wire  _T_11965; // @[StoreQueue.scala 209:52:@7261.6]
  wire  _T_11966; // @[StoreQueue.scala 209:81:@7262.6]
  wire  _T_11969; // @[StoreQueue.scala 209:52:@7264.6]
  wire  _T_11970; // @[StoreQueue.scala 209:81:@7265.6]
  wire  _T_11981; // @[StoreQueue.scala 210:30:@7270.6]
  wire [1:0] _T_11982; // @[OneHot.scala 18:45:@7272.8]
  wire  _T_11983; // @[CircuitMath.scala 30:8:@7273.8]
  wire [31:0] _GEN_1161; // @[StoreQueue.scala 211:30:@7274.8]
  wire [31:0] _GEN_1162; // @[StoreQueue.scala 210:40:@7271.6]
  wire  _GEN_1163; // @[StoreQueue.scala 210:40:@7271.6]
  wire  _T_11988; // @[StoreQueue.scala 215:52:@7278.6]
  wire  _T_11989; // @[StoreQueue.scala 215:81:@7279.6]
  wire  _T_11992; // @[StoreQueue.scala 215:52:@7281.6]
  wire  _T_11993; // @[StoreQueue.scala 215:81:@7282.6]
  wire  _T_12004; // @[StoreQueue.scala 216:30:@7287.6]
  wire [1:0] _T_12005; // @[OneHot.scala 18:45:@7289.8]
  wire  _T_12006; // @[CircuitMath.scala 30:8:@7290.8]
  wire [31:0] _GEN_1165; // @[StoreQueue.scala 217:30:@7291.8]
  wire [31:0] _GEN_1166; // @[StoreQueue.scala 216:40:@7288.6]
  wire  _GEN_1167; // @[StoreQueue.scala 216:40:@7288.6]
  wire  _GEN_1168; // @[StoreQueue.scala 204:35:@7255.4]
  wire  _GEN_1169; // @[StoreQueue.scala 204:35:@7255.4]
  wire [31:0] _GEN_1170; // @[StoreQueue.scala 204:35:@7255.4]
  wire [31:0] _GEN_1171; // @[StoreQueue.scala 204:35:@7255.4]
  wire  _T_12013; // @[StoreQueue.scala 209:52:@7301.6]
  wire  _T_12014; // @[StoreQueue.scala 209:81:@7302.6]
  wire  _T_12017; // @[StoreQueue.scala 209:52:@7304.6]
  wire  _T_12018; // @[StoreQueue.scala 209:81:@7305.6]
  wire  _T_12029; // @[StoreQueue.scala 210:30:@7310.6]
  wire [1:0] _T_12030; // @[OneHot.scala 18:45:@7312.8]
  wire  _T_12031; // @[CircuitMath.scala 30:8:@7313.8]
  wire [31:0] _GEN_1173; // @[StoreQueue.scala 211:30:@7314.8]
  wire [31:0] _GEN_1174; // @[StoreQueue.scala 210:40:@7311.6]
  wire  _GEN_1175; // @[StoreQueue.scala 210:40:@7311.6]
  wire  _T_12036; // @[StoreQueue.scala 215:52:@7318.6]
  wire  _T_12037; // @[StoreQueue.scala 215:81:@7319.6]
  wire  _T_12040; // @[StoreQueue.scala 215:52:@7321.6]
  wire  _T_12041; // @[StoreQueue.scala 215:81:@7322.6]
  wire  _T_12052; // @[StoreQueue.scala 216:30:@7327.6]
  wire [1:0] _T_12053; // @[OneHot.scala 18:45:@7329.8]
  wire  _T_12054; // @[CircuitMath.scala 30:8:@7330.8]
  wire [31:0] _GEN_1177; // @[StoreQueue.scala 217:30:@7331.8]
  wire [31:0] _GEN_1178; // @[StoreQueue.scala 216:40:@7328.6]
  wire  _GEN_1179; // @[StoreQueue.scala 216:40:@7328.6]
  wire  _GEN_1180; // @[StoreQueue.scala 204:35:@7295.4]
  wire  _GEN_1181; // @[StoreQueue.scala 204:35:@7295.4]
  wire [31:0] _GEN_1182; // @[StoreQueue.scala 204:35:@7295.4]
  wire [31:0] _GEN_1183; // @[StoreQueue.scala 204:35:@7295.4]
  wire  _T_12057; // @[StoreQueue.scala 229:23:@7335.4]
  wire [4:0] _T_12060; // @[util.scala 10:8:@7337.6]
  wire [4:0] _GEN_544; // @[util.scala 10:14:@7338.6]
  wire [4:0] _T_12061; // @[util.scala 10:14:@7338.6]
  wire [4:0] _GEN_1184; // @[StoreQueue.scala 229:50:@7336.4]
  wire [3:0] _GEN_1298; // @[util.scala 10:8:@7342.6]
  wire [4:0] _T_12063; // @[util.scala 10:8:@7342.6]
  wire [4:0] _GEN_545; // @[util.scala 10:14:@7343.6]
  wire [4:0] _T_12064; // @[util.scala 10:14:@7343.6]
  wire [4:0] _GEN_1185; // @[StoreQueue.scala 233:20:@7341.4]
  wire  _T_12066; // @[StoreQueue.scala 237:84:@7346.4]
  wire  _T_12067; // @[StoreQueue.scala 237:81:@7347.4]
  wire  _T_12069; // @[StoreQueue.scala 237:84:@7348.4]
  wire  _T_12070; // @[StoreQueue.scala 237:81:@7349.4]
  wire  _T_12072; // @[StoreQueue.scala 237:84:@7350.4]
  wire  _T_12073; // @[StoreQueue.scala 237:81:@7351.4]
  wire  _T_12075; // @[StoreQueue.scala 237:84:@7352.4]
  wire  _T_12076; // @[StoreQueue.scala 237:81:@7353.4]
  wire  _T_12078; // @[StoreQueue.scala 237:84:@7354.4]
  wire  _T_12079; // @[StoreQueue.scala 237:81:@7355.4]
  wire  _T_12081; // @[StoreQueue.scala 237:84:@7356.4]
  wire  _T_12082; // @[StoreQueue.scala 237:81:@7357.4]
  wire  _T_12084; // @[StoreQueue.scala 237:84:@7358.4]
  wire  _T_12085; // @[StoreQueue.scala 237:81:@7359.4]
  wire  _T_12087; // @[StoreQueue.scala 237:84:@7360.4]
  wire  _T_12088; // @[StoreQueue.scala 237:81:@7361.4]
  wire  _T_12090; // @[StoreQueue.scala 237:84:@7362.4]
  wire  _T_12091; // @[StoreQueue.scala 237:81:@7363.4]
  wire  _T_12093; // @[StoreQueue.scala 237:84:@7364.4]
  wire  _T_12094; // @[StoreQueue.scala 237:81:@7365.4]
  wire  _T_12096; // @[StoreQueue.scala 237:84:@7366.4]
  wire  _T_12097; // @[StoreQueue.scala 237:81:@7367.4]
  wire  _T_12099; // @[StoreQueue.scala 237:84:@7368.4]
  wire  _T_12100; // @[StoreQueue.scala 237:81:@7369.4]
  wire  _T_12102; // @[StoreQueue.scala 237:84:@7370.4]
  wire  _T_12103; // @[StoreQueue.scala 237:81:@7371.4]
  wire  _T_12105; // @[StoreQueue.scala 237:84:@7372.4]
  wire  _T_12106; // @[StoreQueue.scala 237:81:@7373.4]
  wire  _T_12108; // @[StoreQueue.scala 237:84:@7374.4]
  wire  _T_12109; // @[StoreQueue.scala 237:81:@7375.4]
  wire  _T_12111; // @[StoreQueue.scala 237:84:@7376.4]
  wire  _T_12112; // @[StoreQueue.scala 237:81:@7377.4]
  wire  _T_12137; // @[StoreQueue.scala 237:98:@7396.4]
  wire  _T_12138; // @[StoreQueue.scala 237:98:@7397.4]
  wire  _T_12139; // @[StoreQueue.scala 237:98:@7398.4]
  wire  _T_12140; // @[StoreQueue.scala 237:98:@7399.4]
  wire  _T_12141; // @[StoreQueue.scala 237:98:@7400.4]
  wire  _T_12142; // @[StoreQueue.scala 237:98:@7401.4]
  wire  _T_12143; // @[StoreQueue.scala 237:98:@7402.4]
  wire  _T_12144; // @[StoreQueue.scala 237:98:@7403.4]
  wire  _T_12145; // @[StoreQueue.scala 237:98:@7404.4]
  wire  _T_12146; // @[StoreQueue.scala 237:98:@7405.4]
  wire  _T_12147; // @[StoreQueue.scala 237:98:@7406.4]
  wire  _T_12148; // @[StoreQueue.scala 237:98:@7407.4]
  wire  _T_12149; // @[StoreQueue.scala 237:98:@7408.4]
  wire  _T_12150; // @[StoreQueue.scala 237:98:@7409.4]
  wire [31:0] _GEN_1187; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1188; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1189; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1190; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1191; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1192; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1193; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1194; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1195; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1196; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1197; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1198; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1199; // @[StoreQueue.scala 252:21:@7479.4]
  wire [31:0] _GEN_1200; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1202 = {{2'd0}, tail}; // @[util.scala 14:20:@173.4]
  assign _T_1604 = 6'h10 - _GEN_1202; // @[util.scala 14:20:@173.4]
  assign _T_1605 = $unsigned(_T_1604); // @[util.scala 14:20:@174.4]
  assign _T_1606 = _T_1605[5:0]; // @[util.scala 14:20:@175.4]
  assign _GEN_0 = _T_1606 % 6'h10; // @[util.scala 14:25:@176.4]
  assign _T_1607 = _GEN_0[4:0]; // @[util.scala 14:25:@176.4]
  assign _GEN_1203 = {{4'd0}, io_bbNumStores}; // @[StoreQueue.scala 70:46:@177.4]
  assign _T_1608 = _T_1607 < _GEN_1203; // @[StoreQueue.scala 70:46:@177.4]
  assign initBits_0 = _T_1608 & io_bbStart; // @[StoreQueue.scala 70:64:@178.4]
  assign _T_1613 = 6'h11 - _GEN_1202; // @[util.scala 14:20:@180.4]
  assign _T_1614 = $unsigned(_T_1613); // @[util.scala 14:20:@181.4]
  assign _T_1615 = _T_1614[5:0]; // @[util.scala 14:20:@182.4]
  assign _GEN_16 = _T_1615 % 6'h10; // @[util.scala 14:25:@183.4]
  assign _T_1616 = _GEN_16[4:0]; // @[util.scala 14:25:@183.4]
  assign _T_1617 = _T_1616 < _GEN_1203; // @[StoreQueue.scala 70:46:@184.4]
  assign initBits_1 = _T_1617 & io_bbStart; // @[StoreQueue.scala 70:64:@185.4]
  assign _T_1622 = 6'h12 - _GEN_1202; // @[util.scala 14:20:@187.4]
  assign _T_1623 = $unsigned(_T_1622); // @[util.scala 14:20:@188.4]
  assign _T_1624 = _T_1623[5:0]; // @[util.scala 14:20:@189.4]
  assign _GEN_34 = _T_1624 % 6'h10; // @[util.scala 14:25:@190.4]
  assign _T_1625 = _GEN_34[4:0]; // @[util.scala 14:25:@190.4]
  assign _T_1626 = _T_1625 < _GEN_1203; // @[StoreQueue.scala 70:46:@191.4]
  assign initBits_2 = _T_1626 & io_bbStart; // @[StoreQueue.scala 70:64:@192.4]
  assign _T_1631 = 6'h13 - _GEN_1202; // @[util.scala 14:20:@194.4]
  assign _T_1632 = $unsigned(_T_1631); // @[util.scala 14:20:@195.4]
  assign _T_1633 = _T_1632[5:0]; // @[util.scala 14:20:@196.4]
  assign _GEN_50 = _T_1633 % 6'h10; // @[util.scala 14:25:@197.4]
  assign _T_1634 = _GEN_50[4:0]; // @[util.scala 14:25:@197.4]
  assign _T_1635 = _T_1634 < _GEN_1203; // @[StoreQueue.scala 70:46:@198.4]
  assign initBits_3 = _T_1635 & io_bbStart; // @[StoreQueue.scala 70:64:@199.4]
  assign _T_1640 = 6'h14 - _GEN_1202; // @[util.scala 14:20:@201.4]
  assign _T_1641 = $unsigned(_T_1640); // @[util.scala 14:20:@202.4]
  assign _T_1642 = _T_1641[5:0]; // @[util.scala 14:20:@203.4]
  assign _GEN_68 = _T_1642 % 6'h10; // @[util.scala 14:25:@204.4]
  assign _T_1643 = _GEN_68[4:0]; // @[util.scala 14:25:@204.4]
  assign _T_1644 = _T_1643 < _GEN_1203; // @[StoreQueue.scala 70:46:@205.4]
  assign initBits_4 = _T_1644 & io_bbStart; // @[StoreQueue.scala 70:64:@206.4]
  assign _T_1649 = 6'h15 - _GEN_1202; // @[util.scala 14:20:@208.4]
  assign _T_1650 = $unsigned(_T_1649); // @[util.scala 14:20:@209.4]
  assign _T_1651 = _T_1650[5:0]; // @[util.scala 14:20:@210.4]
  assign _GEN_84 = _T_1651 % 6'h10; // @[util.scala 14:25:@211.4]
  assign _T_1652 = _GEN_84[4:0]; // @[util.scala 14:25:@211.4]
  assign _T_1653 = _T_1652 < _GEN_1203; // @[StoreQueue.scala 70:46:@212.4]
  assign initBits_5 = _T_1653 & io_bbStart; // @[StoreQueue.scala 70:64:@213.4]
  assign _T_1658 = 6'h16 - _GEN_1202; // @[util.scala 14:20:@215.4]
  assign _T_1659 = $unsigned(_T_1658); // @[util.scala 14:20:@216.4]
  assign _T_1660 = _T_1659[5:0]; // @[util.scala 14:20:@217.4]
  assign _GEN_102 = _T_1660 % 6'h10; // @[util.scala 14:25:@218.4]
  assign _T_1661 = _GEN_102[4:0]; // @[util.scala 14:25:@218.4]
  assign _T_1662 = _T_1661 < _GEN_1203; // @[StoreQueue.scala 70:46:@219.4]
  assign initBits_6 = _T_1662 & io_bbStart; // @[StoreQueue.scala 70:64:@220.4]
  assign _T_1667 = 6'h17 - _GEN_1202; // @[util.scala 14:20:@222.4]
  assign _T_1668 = $unsigned(_T_1667); // @[util.scala 14:20:@223.4]
  assign _T_1669 = _T_1668[5:0]; // @[util.scala 14:20:@224.4]
  assign _GEN_118 = _T_1669 % 6'h10; // @[util.scala 14:25:@225.4]
  assign _T_1670 = _GEN_118[4:0]; // @[util.scala 14:25:@225.4]
  assign _T_1671 = _T_1670 < _GEN_1203; // @[StoreQueue.scala 70:46:@226.4]
  assign initBits_7 = _T_1671 & io_bbStart; // @[StoreQueue.scala 70:64:@227.4]
  assign _T_1676 = 6'h18 - _GEN_1202; // @[util.scala 14:20:@229.4]
  assign _T_1677 = $unsigned(_T_1676); // @[util.scala 14:20:@230.4]
  assign _T_1678 = _T_1677[5:0]; // @[util.scala 14:20:@231.4]
  assign _GEN_136 = _T_1678 % 6'h10; // @[util.scala 14:25:@232.4]
  assign _T_1679 = _GEN_136[4:0]; // @[util.scala 14:25:@232.4]
  assign _T_1680 = _T_1679 < _GEN_1203; // @[StoreQueue.scala 70:46:@233.4]
  assign initBits_8 = _T_1680 & io_bbStart; // @[StoreQueue.scala 70:64:@234.4]
  assign _T_1685 = 6'h19 - _GEN_1202; // @[util.scala 14:20:@236.4]
  assign _T_1686 = $unsigned(_T_1685); // @[util.scala 14:20:@237.4]
  assign _T_1687 = _T_1686[5:0]; // @[util.scala 14:20:@238.4]
  assign _GEN_152 = _T_1687 % 6'h10; // @[util.scala 14:25:@239.4]
  assign _T_1688 = _GEN_152[4:0]; // @[util.scala 14:25:@239.4]
  assign _T_1689 = _T_1688 < _GEN_1203; // @[StoreQueue.scala 70:46:@240.4]
  assign initBits_9 = _T_1689 & io_bbStart; // @[StoreQueue.scala 70:64:@241.4]
  assign _T_1694 = 6'h1a - _GEN_1202; // @[util.scala 14:20:@243.4]
  assign _T_1695 = $unsigned(_T_1694); // @[util.scala 14:20:@244.4]
  assign _T_1696 = _T_1695[5:0]; // @[util.scala 14:20:@245.4]
  assign _GEN_170 = _T_1696 % 6'h10; // @[util.scala 14:25:@246.4]
  assign _T_1697 = _GEN_170[4:0]; // @[util.scala 14:25:@246.4]
  assign _T_1698 = _T_1697 < _GEN_1203; // @[StoreQueue.scala 70:46:@247.4]
  assign initBits_10 = _T_1698 & io_bbStart; // @[StoreQueue.scala 70:64:@248.4]
  assign _T_1703 = 6'h1b - _GEN_1202; // @[util.scala 14:20:@250.4]
  assign _T_1704 = $unsigned(_T_1703); // @[util.scala 14:20:@251.4]
  assign _T_1705 = _T_1704[5:0]; // @[util.scala 14:20:@252.4]
  assign _GEN_186 = _T_1705 % 6'h10; // @[util.scala 14:25:@253.4]
  assign _T_1706 = _GEN_186[4:0]; // @[util.scala 14:25:@253.4]
  assign _T_1707 = _T_1706 < _GEN_1203; // @[StoreQueue.scala 70:46:@254.4]
  assign initBits_11 = _T_1707 & io_bbStart; // @[StoreQueue.scala 70:64:@255.4]
  assign _T_1712 = 6'h1c - _GEN_1202; // @[util.scala 14:20:@257.4]
  assign _T_1713 = $unsigned(_T_1712); // @[util.scala 14:20:@258.4]
  assign _T_1714 = _T_1713[5:0]; // @[util.scala 14:20:@259.4]
  assign _GEN_204 = _T_1714 % 6'h10; // @[util.scala 14:25:@260.4]
  assign _T_1715 = _GEN_204[4:0]; // @[util.scala 14:25:@260.4]
  assign _T_1716 = _T_1715 < _GEN_1203; // @[StoreQueue.scala 70:46:@261.4]
  assign initBits_12 = _T_1716 & io_bbStart; // @[StoreQueue.scala 70:64:@262.4]
  assign _T_1721 = 6'h1d - _GEN_1202; // @[util.scala 14:20:@264.4]
  assign _T_1722 = $unsigned(_T_1721); // @[util.scala 14:20:@265.4]
  assign _T_1723 = _T_1722[5:0]; // @[util.scala 14:20:@266.4]
  assign _GEN_220 = _T_1723 % 6'h10; // @[util.scala 14:25:@267.4]
  assign _T_1724 = _GEN_220[4:0]; // @[util.scala 14:25:@267.4]
  assign _T_1725 = _T_1724 < _GEN_1203; // @[StoreQueue.scala 70:46:@268.4]
  assign initBits_13 = _T_1725 & io_bbStart; // @[StoreQueue.scala 70:64:@269.4]
  assign _T_1730 = 6'h1e - _GEN_1202; // @[util.scala 14:20:@271.4]
  assign _T_1731 = $unsigned(_T_1730); // @[util.scala 14:20:@272.4]
  assign _T_1732 = _T_1731[5:0]; // @[util.scala 14:20:@273.4]
  assign _GEN_238 = _T_1732 % 6'h10; // @[util.scala 14:25:@274.4]
  assign _T_1733 = _GEN_238[4:0]; // @[util.scala 14:25:@274.4]
  assign _T_1734 = _T_1733 < _GEN_1203; // @[StoreQueue.scala 70:46:@275.4]
  assign initBits_14 = _T_1734 & io_bbStart; // @[StoreQueue.scala 70:64:@276.4]
  assign _T_1739 = 6'h1f - _GEN_1202; // @[util.scala 14:20:@278.4]
  assign _T_1740 = $unsigned(_T_1739); // @[util.scala 14:20:@279.4]
  assign _T_1741 = _T_1740[5:0]; // @[util.scala 14:20:@280.4]
  assign _GEN_254 = _T_1741 % 6'h10; // @[util.scala 14:25:@281.4]
  assign _T_1742 = _GEN_254[4:0]; // @[util.scala 14:25:@281.4]
  assign _T_1743 = _T_1742 < _GEN_1203; // @[StoreQueue.scala 70:46:@282.4]
  assign initBits_15 = _T_1743 & io_bbStart; // @[StoreQueue.scala 70:64:@283.4]
  assign _T_1766 = allocatedEntries_0 | initBits_0; // @[StoreQueue.scala 72:78:@301.4]
  assign _T_1767 = allocatedEntries_1 | initBits_1; // @[StoreQueue.scala 72:78:@302.4]
  assign _T_1768 = allocatedEntries_2 | initBits_2; // @[StoreQueue.scala 72:78:@303.4]
  assign _T_1769 = allocatedEntries_3 | initBits_3; // @[StoreQueue.scala 72:78:@304.4]
  assign _T_1770 = allocatedEntries_4 | initBits_4; // @[StoreQueue.scala 72:78:@305.4]
  assign _T_1771 = allocatedEntries_5 | initBits_5; // @[StoreQueue.scala 72:78:@306.4]
  assign _T_1772 = allocatedEntries_6 | initBits_6; // @[StoreQueue.scala 72:78:@307.4]
  assign _T_1773 = allocatedEntries_7 | initBits_7; // @[StoreQueue.scala 72:78:@308.4]
  assign _T_1774 = allocatedEntries_8 | initBits_8; // @[StoreQueue.scala 72:78:@309.4]
  assign _T_1775 = allocatedEntries_9 | initBits_9; // @[StoreQueue.scala 72:78:@310.4]
  assign _T_1776 = allocatedEntries_10 | initBits_10; // @[StoreQueue.scala 72:78:@311.4]
  assign _T_1777 = allocatedEntries_11 | initBits_11; // @[StoreQueue.scala 72:78:@312.4]
  assign _T_1778 = allocatedEntries_12 | initBits_12; // @[StoreQueue.scala 72:78:@313.4]
  assign _T_1779 = allocatedEntries_13 | initBits_13; // @[StoreQueue.scala 72:78:@314.4]
  assign _T_1780 = allocatedEntries_14 | initBits_14; // @[StoreQueue.scala 72:78:@315.4]
  assign _T_1781 = allocatedEntries_15 | initBits_15; // @[StoreQueue.scala 72:78:@316.4]
  assign _T_1812 = _T_1607[3:0]; // @[:@356.6]
  assign _GEN_1 = 4'h1 == _T_1812 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_2 = 4'h2 == _T_1812 ? io_bbStoreOffsets_2 : _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_3 = 4'h3 == _T_1812 ? io_bbStoreOffsets_3 : _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_4 = 4'h4 == _T_1812 ? io_bbStoreOffsets_4 : _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_5 = 4'h5 == _T_1812 ? io_bbStoreOffsets_5 : _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_6 = 4'h6 == _T_1812 ? io_bbStoreOffsets_6 : _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_7 = 4'h7 == _T_1812 ? io_bbStoreOffsets_7 : _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_8 = 4'h8 == _T_1812 ? io_bbStoreOffsets_8 : _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_9 = 4'h9 == _T_1812 ? io_bbStoreOffsets_9 : _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_10 = 4'ha == _T_1812 ? io_bbStoreOffsets_10 : _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_11 = 4'hb == _T_1812 ? io_bbStoreOffsets_11 : _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_12 = 4'hc == _T_1812 ? io_bbStoreOffsets_12 : _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_13 = 4'hd == _T_1812 ? io_bbStoreOffsets_13 : _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_14 = 4'he == _T_1812 ? io_bbStoreOffsets_14 : _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_15 = 4'hf == _T_1812 ? io_bbStoreOffsets_15 : _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_17 = 4'h1 == _T_1812 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_18 = 4'h2 == _T_1812 ? 1'h0 : _GEN_17; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_19 = 4'h3 == _T_1812 ? 1'h0 : _GEN_18; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_20 = 4'h4 == _T_1812 ? 1'h0 : _GEN_19; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_21 = 4'h5 == _T_1812 ? 1'h0 : _GEN_20; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_22 = 4'h6 == _T_1812 ? 1'h0 : _GEN_21; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_23 = 4'h7 == _T_1812 ? 1'h0 : _GEN_22; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_24 = 4'h8 == _T_1812 ? 1'h0 : _GEN_23; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_25 = 4'h9 == _T_1812 ? 1'h0 : _GEN_24; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_26 = 4'ha == _T_1812 ? 1'h0 : _GEN_25; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_27 = 4'hb == _T_1812 ? 1'h0 : _GEN_26; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_28 = 4'hc == _T_1812 ? 1'h0 : _GEN_27; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_29 = 4'hd == _T_1812 ? 1'h0 : _GEN_28; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_30 = 4'he == _T_1812 ? 1'h0 : _GEN_29; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_31 = 4'hf == _T_1812 ? 1'h0 : _GEN_30; // @[StoreQueue.scala 77:18:@364.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _GEN_33 = initBits_0 ? _GEN_31 : portQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _T_1830 = _T_1616[3:0]; // @[:@372.6]
  assign _GEN_35 = 4'h1 == _T_1830 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_36 = 4'h2 == _T_1830 ? io_bbStoreOffsets_2 : _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_37 = 4'h3 == _T_1830 ? io_bbStoreOffsets_3 : _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_38 = 4'h4 == _T_1830 ? io_bbStoreOffsets_4 : _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_39 = 4'h5 == _T_1830 ? io_bbStoreOffsets_5 : _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_40 = 4'h6 == _T_1830 ? io_bbStoreOffsets_6 : _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_41 = 4'h7 == _T_1830 ? io_bbStoreOffsets_7 : _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_42 = 4'h8 == _T_1830 ? io_bbStoreOffsets_8 : _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_43 = 4'h9 == _T_1830 ? io_bbStoreOffsets_9 : _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_44 = 4'ha == _T_1830 ? io_bbStoreOffsets_10 : _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_45 = 4'hb == _T_1830 ? io_bbStoreOffsets_11 : _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_46 = 4'hc == _T_1830 ? io_bbStoreOffsets_12 : _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_47 = 4'hd == _T_1830 ? io_bbStoreOffsets_13 : _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_48 = 4'he == _T_1830 ? io_bbStoreOffsets_14 : _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_49 = 4'hf == _T_1830 ? io_bbStoreOffsets_15 : _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_51 = 4'h1 == _T_1830 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_52 = 4'h2 == _T_1830 ? 1'h0 : _GEN_51; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_53 = 4'h3 == _T_1830 ? 1'h0 : _GEN_52; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_54 = 4'h4 == _T_1830 ? 1'h0 : _GEN_53; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_55 = 4'h5 == _T_1830 ? 1'h0 : _GEN_54; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_56 = 4'h6 == _T_1830 ? 1'h0 : _GEN_55; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_57 = 4'h7 == _T_1830 ? 1'h0 : _GEN_56; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_58 = 4'h8 == _T_1830 ? 1'h0 : _GEN_57; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_59 = 4'h9 == _T_1830 ? 1'h0 : _GEN_58; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_60 = 4'ha == _T_1830 ? 1'h0 : _GEN_59; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_61 = 4'hb == _T_1830 ? 1'h0 : _GEN_60; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_62 = 4'hc == _T_1830 ? 1'h0 : _GEN_61; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_63 = 4'hd == _T_1830 ? 1'h0 : _GEN_62; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_64 = 4'he == _T_1830 ? 1'h0 : _GEN_63; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_65 = 4'hf == _T_1830 ? 1'h0 : _GEN_64; // @[StoreQueue.scala 77:18:@380.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _GEN_67 = initBits_1 ? _GEN_65 : portQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _T_1848 = _T_1625[3:0]; // @[:@388.6]
  assign _GEN_69 = 4'h1 == _T_1848 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_70 = 4'h2 == _T_1848 ? io_bbStoreOffsets_2 : _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_71 = 4'h3 == _T_1848 ? io_bbStoreOffsets_3 : _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_72 = 4'h4 == _T_1848 ? io_bbStoreOffsets_4 : _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_73 = 4'h5 == _T_1848 ? io_bbStoreOffsets_5 : _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_74 = 4'h6 == _T_1848 ? io_bbStoreOffsets_6 : _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_75 = 4'h7 == _T_1848 ? io_bbStoreOffsets_7 : _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_76 = 4'h8 == _T_1848 ? io_bbStoreOffsets_8 : _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_77 = 4'h9 == _T_1848 ? io_bbStoreOffsets_9 : _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_78 = 4'ha == _T_1848 ? io_bbStoreOffsets_10 : _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_79 = 4'hb == _T_1848 ? io_bbStoreOffsets_11 : _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_80 = 4'hc == _T_1848 ? io_bbStoreOffsets_12 : _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_81 = 4'hd == _T_1848 ? io_bbStoreOffsets_13 : _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_82 = 4'he == _T_1848 ? io_bbStoreOffsets_14 : _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_83 = 4'hf == _T_1848 ? io_bbStoreOffsets_15 : _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_85 = 4'h1 == _T_1848 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_86 = 4'h2 == _T_1848 ? 1'h0 : _GEN_85; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_87 = 4'h3 == _T_1848 ? 1'h0 : _GEN_86; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_88 = 4'h4 == _T_1848 ? 1'h0 : _GEN_87; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_89 = 4'h5 == _T_1848 ? 1'h0 : _GEN_88; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_90 = 4'h6 == _T_1848 ? 1'h0 : _GEN_89; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_91 = 4'h7 == _T_1848 ? 1'h0 : _GEN_90; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_92 = 4'h8 == _T_1848 ? 1'h0 : _GEN_91; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_93 = 4'h9 == _T_1848 ? 1'h0 : _GEN_92; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_94 = 4'ha == _T_1848 ? 1'h0 : _GEN_93; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_95 = 4'hb == _T_1848 ? 1'h0 : _GEN_94; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_96 = 4'hc == _T_1848 ? 1'h0 : _GEN_95; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_97 = 4'hd == _T_1848 ? 1'h0 : _GEN_96; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_98 = 4'he == _T_1848 ? 1'h0 : _GEN_97; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_99 = 4'hf == _T_1848 ? 1'h0 : _GEN_98; // @[StoreQueue.scala 77:18:@396.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _GEN_101 = initBits_2 ? _GEN_99 : portQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _T_1866 = _T_1634[3:0]; // @[:@404.6]
  assign _GEN_103 = 4'h1 == _T_1866 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_104 = 4'h2 == _T_1866 ? io_bbStoreOffsets_2 : _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_105 = 4'h3 == _T_1866 ? io_bbStoreOffsets_3 : _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_106 = 4'h4 == _T_1866 ? io_bbStoreOffsets_4 : _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_107 = 4'h5 == _T_1866 ? io_bbStoreOffsets_5 : _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_108 = 4'h6 == _T_1866 ? io_bbStoreOffsets_6 : _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_109 = 4'h7 == _T_1866 ? io_bbStoreOffsets_7 : _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_110 = 4'h8 == _T_1866 ? io_bbStoreOffsets_8 : _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_111 = 4'h9 == _T_1866 ? io_bbStoreOffsets_9 : _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_112 = 4'ha == _T_1866 ? io_bbStoreOffsets_10 : _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_113 = 4'hb == _T_1866 ? io_bbStoreOffsets_11 : _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_114 = 4'hc == _T_1866 ? io_bbStoreOffsets_12 : _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_115 = 4'hd == _T_1866 ? io_bbStoreOffsets_13 : _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_116 = 4'he == _T_1866 ? io_bbStoreOffsets_14 : _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_117 = 4'hf == _T_1866 ? io_bbStoreOffsets_15 : _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_119 = 4'h1 == _T_1866 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_120 = 4'h2 == _T_1866 ? 1'h0 : _GEN_119; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_121 = 4'h3 == _T_1866 ? 1'h0 : _GEN_120; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_122 = 4'h4 == _T_1866 ? 1'h0 : _GEN_121; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_123 = 4'h5 == _T_1866 ? 1'h0 : _GEN_122; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_124 = 4'h6 == _T_1866 ? 1'h0 : _GEN_123; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_125 = 4'h7 == _T_1866 ? 1'h0 : _GEN_124; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_126 = 4'h8 == _T_1866 ? 1'h0 : _GEN_125; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_127 = 4'h9 == _T_1866 ? 1'h0 : _GEN_126; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_128 = 4'ha == _T_1866 ? 1'h0 : _GEN_127; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_129 = 4'hb == _T_1866 ? 1'h0 : _GEN_128; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_130 = 4'hc == _T_1866 ? 1'h0 : _GEN_129; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_131 = 4'hd == _T_1866 ? 1'h0 : _GEN_130; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_132 = 4'he == _T_1866 ? 1'h0 : _GEN_131; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_133 = 4'hf == _T_1866 ? 1'h0 : _GEN_132; // @[StoreQueue.scala 77:18:@412.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _GEN_135 = initBits_3 ? _GEN_133 : portQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _T_1884 = _T_1643[3:0]; // @[:@420.6]
  assign _GEN_137 = 4'h1 == _T_1884 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_138 = 4'h2 == _T_1884 ? io_bbStoreOffsets_2 : _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_139 = 4'h3 == _T_1884 ? io_bbStoreOffsets_3 : _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_140 = 4'h4 == _T_1884 ? io_bbStoreOffsets_4 : _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_141 = 4'h5 == _T_1884 ? io_bbStoreOffsets_5 : _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_142 = 4'h6 == _T_1884 ? io_bbStoreOffsets_6 : _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_143 = 4'h7 == _T_1884 ? io_bbStoreOffsets_7 : _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_144 = 4'h8 == _T_1884 ? io_bbStoreOffsets_8 : _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_145 = 4'h9 == _T_1884 ? io_bbStoreOffsets_9 : _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_146 = 4'ha == _T_1884 ? io_bbStoreOffsets_10 : _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_147 = 4'hb == _T_1884 ? io_bbStoreOffsets_11 : _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_148 = 4'hc == _T_1884 ? io_bbStoreOffsets_12 : _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_149 = 4'hd == _T_1884 ? io_bbStoreOffsets_13 : _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_150 = 4'he == _T_1884 ? io_bbStoreOffsets_14 : _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_151 = 4'hf == _T_1884 ? io_bbStoreOffsets_15 : _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_153 = 4'h1 == _T_1884 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_154 = 4'h2 == _T_1884 ? 1'h0 : _GEN_153; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_155 = 4'h3 == _T_1884 ? 1'h0 : _GEN_154; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_156 = 4'h4 == _T_1884 ? 1'h0 : _GEN_155; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_157 = 4'h5 == _T_1884 ? 1'h0 : _GEN_156; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_158 = 4'h6 == _T_1884 ? 1'h0 : _GEN_157; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_159 = 4'h7 == _T_1884 ? 1'h0 : _GEN_158; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_160 = 4'h8 == _T_1884 ? 1'h0 : _GEN_159; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_161 = 4'h9 == _T_1884 ? 1'h0 : _GEN_160; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_162 = 4'ha == _T_1884 ? 1'h0 : _GEN_161; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_163 = 4'hb == _T_1884 ? 1'h0 : _GEN_162; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_164 = 4'hc == _T_1884 ? 1'h0 : _GEN_163; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_165 = 4'hd == _T_1884 ? 1'h0 : _GEN_164; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_166 = 4'he == _T_1884 ? 1'h0 : _GEN_165; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_167 = 4'hf == _T_1884 ? 1'h0 : _GEN_166; // @[StoreQueue.scala 77:18:@428.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _GEN_169 = initBits_4 ? _GEN_167 : portQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _T_1902 = _T_1652[3:0]; // @[:@436.6]
  assign _GEN_171 = 4'h1 == _T_1902 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_172 = 4'h2 == _T_1902 ? io_bbStoreOffsets_2 : _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_173 = 4'h3 == _T_1902 ? io_bbStoreOffsets_3 : _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_174 = 4'h4 == _T_1902 ? io_bbStoreOffsets_4 : _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_175 = 4'h5 == _T_1902 ? io_bbStoreOffsets_5 : _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_176 = 4'h6 == _T_1902 ? io_bbStoreOffsets_6 : _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_177 = 4'h7 == _T_1902 ? io_bbStoreOffsets_7 : _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_178 = 4'h8 == _T_1902 ? io_bbStoreOffsets_8 : _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_179 = 4'h9 == _T_1902 ? io_bbStoreOffsets_9 : _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_180 = 4'ha == _T_1902 ? io_bbStoreOffsets_10 : _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_181 = 4'hb == _T_1902 ? io_bbStoreOffsets_11 : _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_182 = 4'hc == _T_1902 ? io_bbStoreOffsets_12 : _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_183 = 4'hd == _T_1902 ? io_bbStoreOffsets_13 : _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_184 = 4'he == _T_1902 ? io_bbStoreOffsets_14 : _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_185 = 4'hf == _T_1902 ? io_bbStoreOffsets_15 : _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_187 = 4'h1 == _T_1902 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_188 = 4'h2 == _T_1902 ? 1'h0 : _GEN_187; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_189 = 4'h3 == _T_1902 ? 1'h0 : _GEN_188; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_190 = 4'h4 == _T_1902 ? 1'h0 : _GEN_189; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_191 = 4'h5 == _T_1902 ? 1'h0 : _GEN_190; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_192 = 4'h6 == _T_1902 ? 1'h0 : _GEN_191; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_193 = 4'h7 == _T_1902 ? 1'h0 : _GEN_192; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_194 = 4'h8 == _T_1902 ? 1'h0 : _GEN_193; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_195 = 4'h9 == _T_1902 ? 1'h0 : _GEN_194; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_196 = 4'ha == _T_1902 ? 1'h0 : _GEN_195; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_197 = 4'hb == _T_1902 ? 1'h0 : _GEN_196; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_198 = 4'hc == _T_1902 ? 1'h0 : _GEN_197; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_199 = 4'hd == _T_1902 ? 1'h0 : _GEN_198; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_200 = 4'he == _T_1902 ? 1'h0 : _GEN_199; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_201 = 4'hf == _T_1902 ? 1'h0 : _GEN_200; // @[StoreQueue.scala 77:18:@444.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _GEN_203 = initBits_5 ? _GEN_201 : portQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _T_1920 = _T_1661[3:0]; // @[:@452.6]
  assign _GEN_205 = 4'h1 == _T_1920 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_206 = 4'h2 == _T_1920 ? io_bbStoreOffsets_2 : _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_207 = 4'h3 == _T_1920 ? io_bbStoreOffsets_3 : _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_208 = 4'h4 == _T_1920 ? io_bbStoreOffsets_4 : _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_209 = 4'h5 == _T_1920 ? io_bbStoreOffsets_5 : _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_210 = 4'h6 == _T_1920 ? io_bbStoreOffsets_6 : _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_211 = 4'h7 == _T_1920 ? io_bbStoreOffsets_7 : _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_212 = 4'h8 == _T_1920 ? io_bbStoreOffsets_8 : _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_213 = 4'h9 == _T_1920 ? io_bbStoreOffsets_9 : _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_214 = 4'ha == _T_1920 ? io_bbStoreOffsets_10 : _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_215 = 4'hb == _T_1920 ? io_bbStoreOffsets_11 : _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_216 = 4'hc == _T_1920 ? io_bbStoreOffsets_12 : _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_217 = 4'hd == _T_1920 ? io_bbStoreOffsets_13 : _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_218 = 4'he == _T_1920 ? io_bbStoreOffsets_14 : _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_219 = 4'hf == _T_1920 ? io_bbStoreOffsets_15 : _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_221 = 4'h1 == _T_1920 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_222 = 4'h2 == _T_1920 ? 1'h0 : _GEN_221; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_223 = 4'h3 == _T_1920 ? 1'h0 : _GEN_222; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_224 = 4'h4 == _T_1920 ? 1'h0 : _GEN_223; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_225 = 4'h5 == _T_1920 ? 1'h0 : _GEN_224; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_226 = 4'h6 == _T_1920 ? 1'h0 : _GEN_225; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_227 = 4'h7 == _T_1920 ? 1'h0 : _GEN_226; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_228 = 4'h8 == _T_1920 ? 1'h0 : _GEN_227; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_229 = 4'h9 == _T_1920 ? 1'h0 : _GEN_228; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_230 = 4'ha == _T_1920 ? 1'h0 : _GEN_229; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_231 = 4'hb == _T_1920 ? 1'h0 : _GEN_230; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_232 = 4'hc == _T_1920 ? 1'h0 : _GEN_231; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_233 = 4'hd == _T_1920 ? 1'h0 : _GEN_232; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_234 = 4'he == _T_1920 ? 1'h0 : _GEN_233; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_235 = 4'hf == _T_1920 ? 1'h0 : _GEN_234; // @[StoreQueue.scala 77:18:@460.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _GEN_237 = initBits_6 ? _GEN_235 : portQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _T_1938 = _T_1670[3:0]; // @[:@468.6]
  assign _GEN_239 = 4'h1 == _T_1938 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_240 = 4'h2 == _T_1938 ? io_bbStoreOffsets_2 : _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_241 = 4'h3 == _T_1938 ? io_bbStoreOffsets_3 : _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_242 = 4'h4 == _T_1938 ? io_bbStoreOffsets_4 : _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_243 = 4'h5 == _T_1938 ? io_bbStoreOffsets_5 : _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_244 = 4'h6 == _T_1938 ? io_bbStoreOffsets_6 : _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_245 = 4'h7 == _T_1938 ? io_bbStoreOffsets_7 : _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_246 = 4'h8 == _T_1938 ? io_bbStoreOffsets_8 : _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_247 = 4'h9 == _T_1938 ? io_bbStoreOffsets_9 : _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_248 = 4'ha == _T_1938 ? io_bbStoreOffsets_10 : _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_249 = 4'hb == _T_1938 ? io_bbStoreOffsets_11 : _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_250 = 4'hc == _T_1938 ? io_bbStoreOffsets_12 : _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_251 = 4'hd == _T_1938 ? io_bbStoreOffsets_13 : _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_252 = 4'he == _T_1938 ? io_bbStoreOffsets_14 : _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_253 = 4'hf == _T_1938 ? io_bbStoreOffsets_15 : _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_255 = 4'h1 == _T_1938 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_256 = 4'h2 == _T_1938 ? 1'h0 : _GEN_255; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_257 = 4'h3 == _T_1938 ? 1'h0 : _GEN_256; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_258 = 4'h4 == _T_1938 ? 1'h0 : _GEN_257; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_259 = 4'h5 == _T_1938 ? 1'h0 : _GEN_258; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_260 = 4'h6 == _T_1938 ? 1'h0 : _GEN_259; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_261 = 4'h7 == _T_1938 ? 1'h0 : _GEN_260; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_262 = 4'h8 == _T_1938 ? 1'h0 : _GEN_261; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_263 = 4'h9 == _T_1938 ? 1'h0 : _GEN_262; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_264 = 4'ha == _T_1938 ? 1'h0 : _GEN_263; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_265 = 4'hb == _T_1938 ? 1'h0 : _GEN_264; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_266 = 4'hc == _T_1938 ? 1'h0 : _GEN_265; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_267 = 4'hd == _T_1938 ? 1'h0 : _GEN_266; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_268 = 4'he == _T_1938 ? 1'h0 : _GEN_267; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_269 = 4'hf == _T_1938 ? 1'h0 : _GEN_268; // @[StoreQueue.scala 77:18:@476.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _GEN_271 = initBits_7 ? _GEN_269 : portQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _T_1956 = _T_1679[3:0]; // @[:@484.6]
  assign _GEN_273 = 4'h1 == _T_1956 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_274 = 4'h2 == _T_1956 ? io_bbStoreOffsets_2 : _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_275 = 4'h3 == _T_1956 ? io_bbStoreOffsets_3 : _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_276 = 4'h4 == _T_1956 ? io_bbStoreOffsets_4 : _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_277 = 4'h5 == _T_1956 ? io_bbStoreOffsets_5 : _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_278 = 4'h6 == _T_1956 ? io_bbStoreOffsets_6 : _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_279 = 4'h7 == _T_1956 ? io_bbStoreOffsets_7 : _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_280 = 4'h8 == _T_1956 ? io_bbStoreOffsets_8 : _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_281 = 4'h9 == _T_1956 ? io_bbStoreOffsets_9 : _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_282 = 4'ha == _T_1956 ? io_bbStoreOffsets_10 : _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_283 = 4'hb == _T_1956 ? io_bbStoreOffsets_11 : _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_284 = 4'hc == _T_1956 ? io_bbStoreOffsets_12 : _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_285 = 4'hd == _T_1956 ? io_bbStoreOffsets_13 : _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_286 = 4'he == _T_1956 ? io_bbStoreOffsets_14 : _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_287 = 4'hf == _T_1956 ? io_bbStoreOffsets_15 : _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_289 = 4'h1 == _T_1956 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_290 = 4'h2 == _T_1956 ? 1'h0 : _GEN_289; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_291 = 4'h3 == _T_1956 ? 1'h0 : _GEN_290; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_292 = 4'h4 == _T_1956 ? 1'h0 : _GEN_291; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_293 = 4'h5 == _T_1956 ? 1'h0 : _GEN_292; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_294 = 4'h6 == _T_1956 ? 1'h0 : _GEN_293; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_295 = 4'h7 == _T_1956 ? 1'h0 : _GEN_294; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_296 = 4'h8 == _T_1956 ? 1'h0 : _GEN_295; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_297 = 4'h9 == _T_1956 ? 1'h0 : _GEN_296; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_298 = 4'ha == _T_1956 ? 1'h0 : _GEN_297; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_299 = 4'hb == _T_1956 ? 1'h0 : _GEN_298; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_300 = 4'hc == _T_1956 ? 1'h0 : _GEN_299; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_301 = 4'hd == _T_1956 ? 1'h0 : _GEN_300; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_302 = 4'he == _T_1956 ? 1'h0 : _GEN_301; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_303 = 4'hf == _T_1956 ? 1'h0 : _GEN_302; // @[StoreQueue.scala 77:18:@492.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _GEN_305 = initBits_8 ? _GEN_303 : portQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _T_1974 = _T_1688[3:0]; // @[:@500.6]
  assign _GEN_307 = 4'h1 == _T_1974 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_308 = 4'h2 == _T_1974 ? io_bbStoreOffsets_2 : _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_309 = 4'h3 == _T_1974 ? io_bbStoreOffsets_3 : _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_310 = 4'h4 == _T_1974 ? io_bbStoreOffsets_4 : _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_311 = 4'h5 == _T_1974 ? io_bbStoreOffsets_5 : _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_312 = 4'h6 == _T_1974 ? io_bbStoreOffsets_6 : _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_313 = 4'h7 == _T_1974 ? io_bbStoreOffsets_7 : _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_314 = 4'h8 == _T_1974 ? io_bbStoreOffsets_8 : _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_315 = 4'h9 == _T_1974 ? io_bbStoreOffsets_9 : _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_316 = 4'ha == _T_1974 ? io_bbStoreOffsets_10 : _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_317 = 4'hb == _T_1974 ? io_bbStoreOffsets_11 : _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_318 = 4'hc == _T_1974 ? io_bbStoreOffsets_12 : _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_319 = 4'hd == _T_1974 ? io_bbStoreOffsets_13 : _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_320 = 4'he == _T_1974 ? io_bbStoreOffsets_14 : _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_321 = 4'hf == _T_1974 ? io_bbStoreOffsets_15 : _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_323 = 4'h1 == _T_1974 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_324 = 4'h2 == _T_1974 ? 1'h0 : _GEN_323; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_325 = 4'h3 == _T_1974 ? 1'h0 : _GEN_324; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_326 = 4'h4 == _T_1974 ? 1'h0 : _GEN_325; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_327 = 4'h5 == _T_1974 ? 1'h0 : _GEN_326; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_328 = 4'h6 == _T_1974 ? 1'h0 : _GEN_327; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_329 = 4'h7 == _T_1974 ? 1'h0 : _GEN_328; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_330 = 4'h8 == _T_1974 ? 1'h0 : _GEN_329; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_331 = 4'h9 == _T_1974 ? 1'h0 : _GEN_330; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_332 = 4'ha == _T_1974 ? 1'h0 : _GEN_331; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_333 = 4'hb == _T_1974 ? 1'h0 : _GEN_332; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_334 = 4'hc == _T_1974 ? 1'h0 : _GEN_333; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_335 = 4'hd == _T_1974 ? 1'h0 : _GEN_334; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_336 = 4'he == _T_1974 ? 1'h0 : _GEN_335; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_337 = 4'hf == _T_1974 ? 1'h0 : _GEN_336; // @[StoreQueue.scala 77:18:@508.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _GEN_339 = initBits_9 ? _GEN_337 : portQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _T_1992 = _T_1697[3:0]; // @[:@516.6]
  assign _GEN_341 = 4'h1 == _T_1992 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_342 = 4'h2 == _T_1992 ? io_bbStoreOffsets_2 : _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_343 = 4'h3 == _T_1992 ? io_bbStoreOffsets_3 : _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_344 = 4'h4 == _T_1992 ? io_bbStoreOffsets_4 : _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_345 = 4'h5 == _T_1992 ? io_bbStoreOffsets_5 : _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_346 = 4'h6 == _T_1992 ? io_bbStoreOffsets_6 : _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_347 = 4'h7 == _T_1992 ? io_bbStoreOffsets_7 : _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_348 = 4'h8 == _T_1992 ? io_bbStoreOffsets_8 : _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_349 = 4'h9 == _T_1992 ? io_bbStoreOffsets_9 : _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_350 = 4'ha == _T_1992 ? io_bbStoreOffsets_10 : _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_351 = 4'hb == _T_1992 ? io_bbStoreOffsets_11 : _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_352 = 4'hc == _T_1992 ? io_bbStoreOffsets_12 : _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_353 = 4'hd == _T_1992 ? io_bbStoreOffsets_13 : _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_354 = 4'he == _T_1992 ? io_bbStoreOffsets_14 : _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_355 = 4'hf == _T_1992 ? io_bbStoreOffsets_15 : _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_357 = 4'h1 == _T_1992 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_358 = 4'h2 == _T_1992 ? 1'h0 : _GEN_357; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_359 = 4'h3 == _T_1992 ? 1'h0 : _GEN_358; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_360 = 4'h4 == _T_1992 ? 1'h0 : _GEN_359; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_361 = 4'h5 == _T_1992 ? 1'h0 : _GEN_360; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_362 = 4'h6 == _T_1992 ? 1'h0 : _GEN_361; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_363 = 4'h7 == _T_1992 ? 1'h0 : _GEN_362; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_364 = 4'h8 == _T_1992 ? 1'h0 : _GEN_363; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_365 = 4'h9 == _T_1992 ? 1'h0 : _GEN_364; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_366 = 4'ha == _T_1992 ? 1'h0 : _GEN_365; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_367 = 4'hb == _T_1992 ? 1'h0 : _GEN_366; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_368 = 4'hc == _T_1992 ? 1'h0 : _GEN_367; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_369 = 4'hd == _T_1992 ? 1'h0 : _GEN_368; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_370 = 4'he == _T_1992 ? 1'h0 : _GEN_369; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_371 = 4'hf == _T_1992 ? 1'h0 : _GEN_370; // @[StoreQueue.scala 77:18:@524.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _GEN_373 = initBits_10 ? _GEN_371 : portQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _T_2010 = _T_1706[3:0]; // @[:@532.6]
  assign _GEN_375 = 4'h1 == _T_2010 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_376 = 4'h2 == _T_2010 ? io_bbStoreOffsets_2 : _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_377 = 4'h3 == _T_2010 ? io_bbStoreOffsets_3 : _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_378 = 4'h4 == _T_2010 ? io_bbStoreOffsets_4 : _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_379 = 4'h5 == _T_2010 ? io_bbStoreOffsets_5 : _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_380 = 4'h6 == _T_2010 ? io_bbStoreOffsets_6 : _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_381 = 4'h7 == _T_2010 ? io_bbStoreOffsets_7 : _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_382 = 4'h8 == _T_2010 ? io_bbStoreOffsets_8 : _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_383 = 4'h9 == _T_2010 ? io_bbStoreOffsets_9 : _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_384 = 4'ha == _T_2010 ? io_bbStoreOffsets_10 : _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_385 = 4'hb == _T_2010 ? io_bbStoreOffsets_11 : _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_386 = 4'hc == _T_2010 ? io_bbStoreOffsets_12 : _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_387 = 4'hd == _T_2010 ? io_bbStoreOffsets_13 : _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_388 = 4'he == _T_2010 ? io_bbStoreOffsets_14 : _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_389 = 4'hf == _T_2010 ? io_bbStoreOffsets_15 : _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_391 = 4'h1 == _T_2010 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_392 = 4'h2 == _T_2010 ? 1'h0 : _GEN_391; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_393 = 4'h3 == _T_2010 ? 1'h0 : _GEN_392; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_394 = 4'h4 == _T_2010 ? 1'h0 : _GEN_393; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_395 = 4'h5 == _T_2010 ? 1'h0 : _GEN_394; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_396 = 4'h6 == _T_2010 ? 1'h0 : _GEN_395; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_397 = 4'h7 == _T_2010 ? 1'h0 : _GEN_396; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_398 = 4'h8 == _T_2010 ? 1'h0 : _GEN_397; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_399 = 4'h9 == _T_2010 ? 1'h0 : _GEN_398; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_400 = 4'ha == _T_2010 ? 1'h0 : _GEN_399; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_401 = 4'hb == _T_2010 ? 1'h0 : _GEN_400; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_402 = 4'hc == _T_2010 ? 1'h0 : _GEN_401; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_403 = 4'hd == _T_2010 ? 1'h0 : _GEN_402; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_404 = 4'he == _T_2010 ? 1'h0 : _GEN_403; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_405 = 4'hf == _T_2010 ? 1'h0 : _GEN_404; // @[StoreQueue.scala 77:18:@540.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _GEN_407 = initBits_11 ? _GEN_405 : portQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _T_2028 = _T_1715[3:0]; // @[:@548.6]
  assign _GEN_409 = 4'h1 == _T_2028 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_410 = 4'h2 == _T_2028 ? io_bbStoreOffsets_2 : _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_411 = 4'h3 == _T_2028 ? io_bbStoreOffsets_3 : _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_412 = 4'h4 == _T_2028 ? io_bbStoreOffsets_4 : _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_413 = 4'h5 == _T_2028 ? io_bbStoreOffsets_5 : _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_414 = 4'h6 == _T_2028 ? io_bbStoreOffsets_6 : _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_415 = 4'h7 == _T_2028 ? io_bbStoreOffsets_7 : _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_416 = 4'h8 == _T_2028 ? io_bbStoreOffsets_8 : _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_417 = 4'h9 == _T_2028 ? io_bbStoreOffsets_9 : _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_418 = 4'ha == _T_2028 ? io_bbStoreOffsets_10 : _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_419 = 4'hb == _T_2028 ? io_bbStoreOffsets_11 : _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_420 = 4'hc == _T_2028 ? io_bbStoreOffsets_12 : _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_421 = 4'hd == _T_2028 ? io_bbStoreOffsets_13 : _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_422 = 4'he == _T_2028 ? io_bbStoreOffsets_14 : _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_423 = 4'hf == _T_2028 ? io_bbStoreOffsets_15 : _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_425 = 4'h1 == _T_2028 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_426 = 4'h2 == _T_2028 ? 1'h0 : _GEN_425; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_427 = 4'h3 == _T_2028 ? 1'h0 : _GEN_426; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_428 = 4'h4 == _T_2028 ? 1'h0 : _GEN_427; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_429 = 4'h5 == _T_2028 ? 1'h0 : _GEN_428; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_430 = 4'h6 == _T_2028 ? 1'h0 : _GEN_429; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_431 = 4'h7 == _T_2028 ? 1'h0 : _GEN_430; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_432 = 4'h8 == _T_2028 ? 1'h0 : _GEN_431; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_433 = 4'h9 == _T_2028 ? 1'h0 : _GEN_432; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_434 = 4'ha == _T_2028 ? 1'h0 : _GEN_433; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_435 = 4'hb == _T_2028 ? 1'h0 : _GEN_434; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_436 = 4'hc == _T_2028 ? 1'h0 : _GEN_435; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_437 = 4'hd == _T_2028 ? 1'h0 : _GEN_436; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_438 = 4'he == _T_2028 ? 1'h0 : _GEN_437; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_439 = 4'hf == _T_2028 ? 1'h0 : _GEN_438; // @[StoreQueue.scala 77:18:@556.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _GEN_441 = initBits_12 ? _GEN_439 : portQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _T_2046 = _T_1724[3:0]; // @[:@564.6]
  assign _GEN_443 = 4'h1 == _T_2046 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_444 = 4'h2 == _T_2046 ? io_bbStoreOffsets_2 : _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_445 = 4'h3 == _T_2046 ? io_bbStoreOffsets_3 : _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_446 = 4'h4 == _T_2046 ? io_bbStoreOffsets_4 : _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_447 = 4'h5 == _T_2046 ? io_bbStoreOffsets_5 : _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_448 = 4'h6 == _T_2046 ? io_bbStoreOffsets_6 : _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_449 = 4'h7 == _T_2046 ? io_bbStoreOffsets_7 : _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_450 = 4'h8 == _T_2046 ? io_bbStoreOffsets_8 : _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_451 = 4'h9 == _T_2046 ? io_bbStoreOffsets_9 : _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_452 = 4'ha == _T_2046 ? io_bbStoreOffsets_10 : _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_453 = 4'hb == _T_2046 ? io_bbStoreOffsets_11 : _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_454 = 4'hc == _T_2046 ? io_bbStoreOffsets_12 : _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_455 = 4'hd == _T_2046 ? io_bbStoreOffsets_13 : _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_456 = 4'he == _T_2046 ? io_bbStoreOffsets_14 : _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_457 = 4'hf == _T_2046 ? io_bbStoreOffsets_15 : _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_459 = 4'h1 == _T_2046 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_460 = 4'h2 == _T_2046 ? 1'h0 : _GEN_459; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_461 = 4'h3 == _T_2046 ? 1'h0 : _GEN_460; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_462 = 4'h4 == _T_2046 ? 1'h0 : _GEN_461; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_463 = 4'h5 == _T_2046 ? 1'h0 : _GEN_462; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_464 = 4'h6 == _T_2046 ? 1'h0 : _GEN_463; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_465 = 4'h7 == _T_2046 ? 1'h0 : _GEN_464; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_466 = 4'h8 == _T_2046 ? 1'h0 : _GEN_465; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_467 = 4'h9 == _T_2046 ? 1'h0 : _GEN_466; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_468 = 4'ha == _T_2046 ? 1'h0 : _GEN_467; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_469 = 4'hb == _T_2046 ? 1'h0 : _GEN_468; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_470 = 4'hc == _T_2046 ? 1'h0 : _GEN_469; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_471 = 4'hd == _T_2046 ? 1'h0 : _GEN_470; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_472 = 4'he == _T_2046 ? 1'h0 : _GEN_471; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_473 = 4'hf == _T_2046 ? 1'h0 : _GEN_472; // @[StoreQueue.scala 77:18:@572.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _GEN_475 = initBits_13 ? _GEN_473 : portQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _T_2064 = _T_1733[3:0]; // @[:@580.6]
  assign _GEN_477 = 4'h1 == _T_2064 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_478 = 4'h2 == _T_2064 ? io_bbStoreOffsets_2 : _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_479 = 4'h3 == _T_2064 ? io_bbStoreOffsets_3 : _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_480 = 4'h4 == _T_2064 ? io_bbStoreOffsets_4 : _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_481 = 4'h5 == _T_2064 ? io_bbStoreOffsets_5 : _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_482 = 4'h6 == _T_2064 ? io_bbStoreOffsets_6 : _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_483 = 4'h7 == _T_2064 ? io_bbStoreOffsets_7 : _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_484 = 4'h8 == _T_2064 ? io_bbStoreOffsets_8 : _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_485 = 4'h9 == _T_2064 ? io_bbStoreOffsets_9 : _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_486 = 4'ha == _T_2064 ? io_bbStoreOffsets_10 : _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_487 = 4'hb == _T_2064 ? io_bbStoreOffsets_11 : _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_488 = 4'hc == _T_2064 ? io_bbStoreOffsets_12 : _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_489 = 4'hd == _T_2064 ? io_bbStoreOffsets_13 : _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_490 = 4'he == _T_2064 ? io_bbStoreOffsets_14 : _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_491 = 4'hf == _T_2064 ? io_bbStoreOffsets_15 : _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_493 = 4'h1 == _T_2064 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_494 = 4'h2 == _T_2064 ? 1'h0 : _GEN_493; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_495 = 4'h3 == _T_2064 ? 1'h0 : _GEN_494; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_496 = 4'h4 == _T_2064 ? 1'h0 : _GEN_495; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_497 = 4'h5 == _T_2064 ? 1'h0 : _GEN_496; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_498 = 4'h6 == _T_2064 ? 1'h0 : _GEN_497; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_499 = 4'h7 == _T_2064 ? 1'h0 : _GEN_498; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_500 = 4'h8 == _T_2064 ? 1'h0 : _GEN_499; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_501 = 4'h9 == _T_2064 ? 1'h0 : _GEN_500; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_502 = 4'ha == _T_2064 ? 1'h0 : _GEN_501; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_503 = 4'hb == _T_2064 ? 1'h0 : _GEN_502; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_504 = 4'hc == _T_2064 ? 1'h0 : _GEN_503; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_505 = 4'hd == _T_2064 ? 1'h0 : _GEN_504; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_506 = 4'he == _T_2064 ? 1'h0 : _GEN_505; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_507 = 4'hf == _T_2064 ? 1'h0 : _GEN_506; // @[StoreQueue.scala 77:18:@588.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _GEN_509 = initBits_14 ? _GEN_507 : portQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _T_2082 = _T_1742[3:0]; // @[:@596.6]
  assign _GEN_511 = 4'h1 == _T_2082 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_512 = 4'h2 == _T_2082 ? io_bbStoreOffsets_2 : _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_513 = 4'h3 == _T_2082 ? io_bbStoreOffsets_3 : _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_514 = 4'h4 == _T_2082 ? io_bbStoreOffsets_4 : _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_515 = 4'h5 == _T_2082 ? io_bbStoreOffsets_5 : _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_516 = 4'h6 == _T_2082 ? io_bbStoreOffsets_6 : _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_517 = 4'h7 == _T_2082 ? io_bbStoreOffsets_7 : _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_518 = 4'h8 == _T_2082 ? io_bbStoreOffsets_8 : _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_519 = 4'h9 == _T_2082 ? io_bbStoreOffsets_9 : _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_520 = 4'ha == _T_2082 ? io_bbStoreOffsets_10 : _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_521 = 4'hb == _T_2082 ? io_bbStoreOffsets_11 : _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_522 = 4'hc == _T_2082 ? io_bbStoreOffsets_12 : _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_523 = 4'hd == _T_2082 ? io_bbStoreOffsets_13 : _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_524 = 4'he == _T_2082 ? io_bbStoreOffsets_14 : _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_525 = 4'hf == _T_2082 ? io_bbStoreOffsets_15 : _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_527 = 4'h1 == _T_2082 ? 1'h0 : io_bbStorePorts_0; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_528 = 4'h2 == _T_2082 ? 1'h0 : _GEN_527; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_529 = 4'h3 == _T_2082 ? 1'h0 : _GEN_528; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_530 = 4'h4 == _T_2082 ? 1'h0 : _GEN_529; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_531 = 4'h5 == _T_2082 ? 1'h0 : _GEN_530; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_532 = 4'h6 == _T_2082 ? 1'h0 : _GEN_531; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_533 = 4'h7 == _T_2082 ? 1'h0 : _GEN_532; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_534 = 4'h8 == _T_2082 ? 1'h0 : _GEN_533; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_535 = 4'h9 == _T_2082 ? 1'h0 : _GEN_534; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_536 = 4'ha == _T_2082 ? 1'h0 : _GEN_535; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_537 = 4'hb == _T_2082 ? 1'h0 : _GEN_536; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_538 = 4'hc == _T_2082 ? 1'h0 : _GEN_537; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_539 = 4'hd == _T_2082 ? 1'h0 : _GEN_538; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_540 = 4'he == _T_2082 ? 1'h0 : _GEN_539; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_541 = 4'hf == _T_2082 ? 1'h0 : _GEN_540; // @[StoreQueue.scala 77:18:@604.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _GEN_543 = initBits_15 ? _GEN_541 : portQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _T_2104 = _GEN_15 + 4'h1; // @[util.scala 10:8:@615.6]
  assign _GEN_272 = _T_2104 % 5'h10; // @[util.scala 10:14:@616.6]
  assign _T_2105 = _GEN_272[4:0]; // @[util.scala 10:14:@616.6]
  assign _GEN_1267 = {{1'd0}, io_loadTail}; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2106 = _T_2105 == _GEN_1267; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2107 = io_loadEmpty & _T_2106; // @[StoreQueue.scala 95:50:@618.6]
  assign _T_2109 = _T_2107 == 1'h0; // @[StoreQueue.scala 95:35:@619.6]
  assign _T_2111 = previousLoadHead <= offsetQ_0; // @[StoreQueue.scala 100:35:@627.8]
  assign _T_2112 = offsetQ_0 < io_loadHead; // @[StoreQueue.scala 100:87:@628.8]
  assign _T_2113 = _T_2111 & _T_2112; // @[StoreQueue.scala 100:61:@629.8]
  assign _T_2115 = previousLoadHead > io_loadHead; // @[StoreQueue.scala 102:35:@634.10]
  assign _T_2116 = io_loadHead <= offsetQ_0; // @[StoreQueue.scala 103:23:@635.10]
  assign _T_2117 = offsetQ_0 < previousLoadHead; // @[StoreQueue.scala 103:75:@636.10]
  assign _T_2118 = _T_2116 & _T_2117; // @[StoreQueue.scala 103:49:@637.10]
  assign _T_2120 = _T_2118 == 1'h0; // @[StoreQueue.scala 103:9:@638.10]
  assign _T_2121 = _T_2115 & _T_2120; // @[StoreQueue.scala 102:49:@639.10]
  assign _GEN_560 = _T_2121 ? 1'h0 : checkBits_0; // @[StoreQueue.scala 103:96:@640.10]
  assign _GEN_561 = _T_2113 ? 1'h0 : _GEN_560; // @[StoreQueue.scala 100:102:@630.8]
  assign _GEN_562 = io_loadEmpty ? 1'h0 : _GEN_561; // @[StoreQueue.scala 98:26:@623.6]
  assign _GEN_563 = initBits_0 ? _T_2109 : _GEN_562; // @[StoreQueue.scala 94:35:@608.4]
  assign _T_2134 = _GEN_49 + 4'h1; // @[util.scala 10:8:@651.6]
  assign _GEN_288 = _T_2134 % 5'h10; // @[util.scala 10:14:@652.6]
  assign _T_2135 = _GEN_288[4:0]; // @[util.scala 10:14:@652.6]
  assign _T_2136 = _T_2135 == _GEN_1267; // @[StoreQueue.scala 96:56:@653.6]
  assign _T_2137 = io_loadEmpty & _T_2136; // @[StoreQueue.scala 95:50:@654.6]
  assign _T_2139 = _T_2137 == 1'h0; // @[StoreQueue.scala 95:35:@655.6]
  assign _T_2141 = previousLoadHead <= offsetQ_1; // @[StoreQueue.scala 100:35:@663.8]
  assign _T_2142 = offsetQ_1 < io_loadHead; // @[StoreQueue.scala 100:87:@664.8]
  assign _T_2143 = _T_2141 & _T_2142; // @[StoreQueue.scala 100:61:@665.8]
  assign _T_2146 = io_loadHead <= offsetQ_1; // @[StoreQueue.scala 103:23:@671.10]
  assign _T_2147 = offsetQ_1 < previousLoadHead; // @[StoreQueue.scala 103:75:@672.10]
  assign _T_2148 = _T_2146 & _T_2147; // @[StoreQueue.scala 103:49:@673.10]
  assign _T_2150 = _T_2148 == 1'h0; // @[StoreQueue.scala 103:9:@674.10]
  assign _T_2151 = _T_2115 & _T_2150; // @[StoreQueue.scala 102:49:@675.10]
  assign _GEN_580 = _T_2151 ? 1'h0 : checkBits_1; // @[StoreQueue.scala 103:96:@676.10]
  assign _GEN_581 = _T_2143 ? 1'h0 : _GEN_580; // @[StoreQueue.scala 100:102:@666.8]
  assign _GEN_582 = io_loadEmpty ? 1'h0 : _GEN_581; // @[StoreQueue.scala 98:26:@659.6]
  assign _GEN_583 = initBits_1 ? _T_2139 : _GEN_582; // @[StoreQueue.scala 94:35:@644.4]
  assign _T_2164 = _GEN_83 + 4'h1; // @[util.scala 10:8:@687.6]
  assign _GEN_306 = _T_2164 % 5'h10; // @[util.scala 10:14:@688.6]
  assign _T_2165 = _GEN_306[4:0]; // @[util.scala 10:14:@688.6]
  assign _T_2166 = _T_2165 == _GEN_1267; // @[StoreQueue.scala 96:56:@689.6]
  assign _T_2167 = io_loadEmpty & _T_2166; // @[StoreQueue.scala 95:50:@690.6]
  assign _T_2169 = _T_2167 == 1'h0; // @[StoreQueue.scala 95:35:@691.6]
  assign _T_2171 = previousLoadHead <= offsetQ_2; // @[StoreQueue.scala 100:35:@699.8]
  assign _T_2172 = offsetQ_2 < io_loadHead; // @[StoreQueue.scala 100:87:@700.8]
  assign _T_2173 = _T_2171 & _T_2172; // @[StoreQueue.scala 100:61:@701.8]
  assign _T_2176 = io_loadHead <= offsetQ_2; // @[StoreQueue.scala 103:23:@707.10]
  assign _T_2177 = offsetQ_2 < previousLoadHead; // @[StoreQueue.scala 103:75:@708.10]
  assign _T_2178 = _T_2176 & _T_2177; // @[StoreQueue.scala 103:49:@709.10]
  assign _T_2180 = _T_2178 == 1'h0; // @[StoreQueue.scala 103:9:@710.10]
  assign _T_2181 = _T_2115 & _T_2180; // @[StoreQueue.scala 102:49:@711.10]
  assign _GEN_600 = _T_2181 ? 1'h0 : checkBits_2; // @[StoreQueue.scala 103:96:@712.10]
  assign _GEN_601 = _T_2173 ? 1'h0 : _GEN_600; // @[StoreQueue.scala 100:102:@702.8]
  assign _GEN_602 = io_loadEmpty ? 1'h0 : _GEN_601; // @[StoreQueue.scala 98:26:@695.6]
  assign _GEN_603 = initBits_2 ? _T_2169 : _GEN_602; // @[StoreQueue.scala 94:35:@680.4]
  assign _T_2194 = _GEN_117 + 4'h1; // @[util.scala 10:8:@723.6]
  assign _GEN_322 = _T_2194 % 5'h10; // @[util.scala 10:14:@724.6]
  assign _T_2195 = _GEN_322[4:0]; // @[util.scala 10:14:@724.6]
  assign _T_2196 = _T_2195 == _GEN_1267; // @[StoreQueue.scala 96:56:@725.6]
  assign _T_2197 = io_loadEmpty & _T_2196; // @[StoreQueue.scala 95:50:@726.6]
  assign _T_2199 = _T_2197 == 1'h0; // @[StoreQueue.scala 95:35:@727.6]
  assign _T_2201 = previousLoadHead <= offsetQ_3; // @[StoreQueue.scala 100:35:@735.8]
  assign _T_2202 = offsetQ_3 < io_loadHead; // @[StoreQueue.scala 100:87:@736.8]
  assign _T_2203 = _T_2201 & _T_2202; // @[StoreQueue.scala 100:61:@737.8]
  assign _T_2206 = io_loadHead <= offsetQ_3; // @[StoreQueue.scala 103:23:@743.10]
  assign _T_2207 = offsetQ_3 < previousLoadHead; // @[StoreQueue.scala 103:75:@744.10]
  assign _T_2208 = _T_2206 & _T_2207; // @[StoreQueue.scala 103:49:@745.10]
  assign _T_2210 = _T_2208 == 1'h0; // @[StoreQueue.scala 103:9:@746.10]
  assign _T_2211 = _T_2115 & _T_2210; // @[StoreQueue.scala 102:49:@747.10]
  assign _GEN_620 = _T_2211 ? 1'h0 : checkBits_3; // @[StoreQueue.scala 103:96:@748.10]
  assign _GEN_621 = _T_2203 ? 1'h0 : _GEN_620; // @[StoreQueue.scala 100:102:@738.8]
  assign _GEN_622 = io_loadEmpty ? 1'h0 : _GEN_621; // @[StoreQueue.scala 98:26:@731.6]
  assign _GEN_623 = initBits_3 ? _T_2199 : _GEN_622; // @[StoreQueue.scala 94:35:@716.4]
  assign _T_2224 = _GEN_151 + 4'h1; // @[util.scala 10:8:@759.6]
  assign _GEN_340 = _T_2224 % 5'h10; // @[util.scala 10:14:@760.6]
  assign _T_2225 = _GEN_340[4:0]; // @[util.scala 10:14:@760.6]
  assign _T_2226 = _T_2225 == _GEN_1267; // @[StoreQueue.scala 96:56:@761.6]
  assign _T_2227 = io_loadEmpty & _T_2226; // @[StoreQueue.scala 95:50:@762.6]
  assign _T_2229 = _T_2227 == 1'h0; // @[StoreQueue.scala 95:35:@763.6]
  assign _T_2231 = previousLoadHead <= offsetQ_4; // @[StoreQueue.scala 100:35:@771.8]
  assign _T_2232 = offsetQ_4 < io_loadHead; // @[StoreQueue.scala 100:87:@772.8]
  assign _T_2233 = _T_2231 & _T_2232; // @[StoreQueue.scala 100:61:@773.8]
  assign _T_2236 = io_loadHead <= offsetQ_4; // @[StoreQueue.scala 103:23:@779.10]
  assign _T_2237 = offsetQ_4 < previousLoadHead; // @[StoreQueue.scala 103:75:@780.10]
  assign _T_2238 = _T_2236 & _T_2237; // @[StoreQueue.scala 103:49:@781.10]
  assign _T_2240 = _T_2238 == 1'h0; // @[StoreQueue.scala 103:9:@782.10]
  assign _T_2241 = _T_2115 & _T_2240; // @[StoreQueue.scala 102:49:@783.10]
  assign _GEN_640 = _T_2241 ? 1'h0 : checkBits_4; // @[StoreQueue.scala 103:96:@784.10]
  assign _GEN_641 = _T_2233 ? 1'h0 : _GEN_640; // @[StoreQueue.scala 100:102:@774.8]
  assign _GEN_642 = io_loadEmpty ? 1'h0 : _GEN_641; // @[StoreQueue.scala 98:26:@767.6]
  assign _GEN_643 = initBits_4 ? _T_2229 : _GEN_642; // @[StoreQueue.scala 94:35:@752.4]
  assign _T_2254 = _GEN_185 + 4'h1; // @[util.scala 10:8:@795.6]
  assign _GEN_356 = _T_2254 % 5'h10; // @[util.scala 10:14:@796.6]
  assign _T_2255 = _GEN_356[4:0]; // @[util.scala 10:14:@796.6]
  assign _T_2256 = _T_2255 == _GEN_1267; // @[StoreQueue.scala 96:56:@797.6]
  assign _T_2257 = io_loadEmpty & _T_2256; // @[StoreQueue.scala 95:50:@798.6]
  assign _T_2259 = _T_2257 == 1'h0; // @[StoreQueue.scala 95:35:@799.6]
  assign _T_2261 = previousLoadHead <= offsetQ_5; // @[StoreQueue.scala 100:35:@807.8]
  assign _T_2262 = offsetQ_5 < io_loadHead; // @[StoreQueue.scala 100:87:@808.8]
  assign _T_2263 = _T_2261 & _T_2262; // @[StoreQueue.scala 100:61:@809.8]
  assign _T_2266 = io_loadHead <= offsetQ_5; // @[StoreQueue.scala 103:23:@815.10]
  assign _T_2267 = offsetQ_5 < previousLoadHead; // @[StoreQueue.scala 103:75:@816.10]
  assign _T_2268 = _T_2266 & _T_2267; // @[StoreQueue.scala 103:49:@817.10]
  assign _T_2270 = _T_2268 == 1'h0; // @[StoreQueue.scala 103:9:@818.10]
  assign _T_2271 = _T_2115 & _T_2270; // @[StoreQueue.scala 102:49:@819.10]
  assign _GEN_660 = _T_2271 ? 1'h0 : checkBits_5; // @[StoreQueue.scala 103:96:@820.10]
  assign _GEN_661 = _T_2263 ? 1'h0 : _GEN_660; // @[StoreQueue.scala 100:102:@810.8]
  assign _GEN_662 = io_loadEmpty ? 1'h0 : _GEN_661; // @[StoreQueue.scala 98:26:@803.6]
  assign _GEN_663 = initBits_5 ? _T_2259 : _GEN_662; // @[StoreQueue.scala 94:35:@788.4]
  assign _T_2284 = _GEN_219 + 4'h1; // @[util.scala 10:8:@831.6]
  assign _GEN_374 = _T_2284 % 5'h10; // @[util.scala 10:14:@832.6]
  assign _T_2285 = _GEN_374[4:0]; // @[util.scala 10:14:@832.6]
  assign _T_2286 = _T_2285 == _GEN_1267; // @[StoreQueue.scala 96:56:@833.6]
  assign _T_2287 = io_loadEmpty & _T_2286; // @[StoreQueue.scala 95:50:@834.6]
  assign _T_2289 = _T_2287 == 1'h0; // @[StoreQueue.scala 95:35:@835.6]
  assign _T_2291 = previousLoadHead <= offsetQ_6; // @[StoreQueue.scala 100:35:@843.8]
  assign _T_2292 = offsetQ_6 < io_loadHead; // @[StoreQueue.scala 100:87:@844.8]
  assign _T_2293 = _T_2291 & _T_2292; // @[StoreQueue.scala 100:61:@845.8]
  assign _T_2296 = io_loadHead <= offsetQ_6; // @[StoreQueue.scala 103:23:@851.10]
  assign _T_2297 = offsetQ_6 < previousLoadHead; // @[StoreQueue.scala 103:75:@852.10]
  assign _T_2298 = _T_2296 & _T_2297; // @[StoreQueue.scala 103:49:@853.10]
  assign _T_2300 = _T_2298 == 1'h0; // @[StoreQueue.scala 103:9:@854.10]
  assign _T_2301 = _T_2115 & _T_2300; // @[StoreQueue.scala 102:49:@855.10]
  assign _GEN_680 = _T_2301 ? 1'h0 : checkBits_6; // @[StoreQueue.scala 103:96:@856.10]
  assign _GEN_681 = _T_2293 ? 1'h0 : _GEN_680; // @[StoreQueue.scala 100:102:@846.8]
  assign _GEN_682 = io_loadEmpty ? 1'h0 : _GEN_681; // @[StoreQueue.scala 98:26:@839.6]
  assign _GEN_683 = initBits_6 ? _T_2289 : _GEN_682; // @[StoreQueue.scala 94:35:@824.4]
  assign _T_2314 = _GEN_253 + 4'h1; // @[util.scala 10:8:@867.6]
  assign _GEN_390 = _T_2314 % 5'h10; // @[util.scala 10:14:@868.6]
  assign _T_2315 = _GEN_390[4:0]; // @[util.scala 10:14:@868.6]
  assign _T_2316 = _T_2315 == _GEN_1267; // @[StoreQueue.scala 96:56:@869.6]
  assign _T_2317 = io_loadEmpty & _T_2316; // @[StoreQueue.scala 95:50:@870.6]
  assign _T_2319 = _T_2317 == 1'h0; // @[StoreQueue.scala 95:35:@871.6]
  assign _T_2321 = previousLoadHead <= offsetQ_7; // @[StoreQueue.scala 100:35:@879.8]
  assign _T_2322 = offsetQ_7 < io_loadHead; // @[StoreQueue.scala 100:87:@880.8]
  assign _T_2323 = _T_2321 & _T_2322; // @[StoreQueue.scala 100:61:@881.8]
  assign _T_2326 = io_loadHead <= offsetQ_7; // @[StoreQueue.scala 103:23:@887.10]
  assign _T_2327 = offsetQ_7 < previousLoadHead; // @[StoreQueue.scala 103:75:@888.10]
  assign _T_2328 = _T_2326 & _T_2327; // @[StoreQueue.scala 103:49:@889.10]
  assign _T_2330 = _T_2328 == 1'h0; // @[StoreQueue.scala 103:9:@890.10]
  assign _T_2331 = _T_2115 & _T_2330; // @[StoreQueue.scala 102:49:@891.10]
  assign _GEN_700 = _T_2331 ? 1'h0 : checkBits_7; // @[StoreQueue.scala 103:96:@892.10]
  assign _GEN_701 = _T_2323 ? 1'h0 : _GEN_700; // @[StoreQueue.scala 100:102:@882.8]
  assign _GEN_702 = io_loadEmpty ? 1'h0 : _GEN_701; // @[StoreQueue.scala 98:26:@875.6]
  assign _GEN_703 = initBits_7 ? _T_2319 : _GEN_702; // @[StoreQueue.scala 94:35:@860.4]
  assign _T_2344 = _GEN_287 + 4'h1; // @[util.scala 10:8:@903.6]
  assign _GEN_408 = _T_2344 % 5'h10; // @[util.scala 10:14:@904.6]
  assign _T_2345 = _GEN_408[4:0]; // @[util.scala 10:14:@904.6]
  assign _T_2346 = _T_2345 == _GEN_1267; // @[StoreQueue.scala 96:56:@905.6]
  assign _T_2347 = io_loadEmpty & _T_2346; // @[StoreQueue.scala 95:50:@906.6]
  assign _T_2349 = _T_2347 == 1'h0; // @[StoreQueue.scala 95:35:@907.6]
  assign _T_2351 = previousLoadHead <= offsetQ_8; // @[StoreQueue.scala 100:35:@915.8]
  assign _T_2352 = offsetQ_8 < io_loadHead; // @[StoreQueue.scala 100:87:@916.8]
  assign _T_2353 = _T_2351 & _T_2352; // @[StoreQueue.scala 100:61:@917.8]
  assign _T_2356 = io_loadHead <= offsetQ_8; // @[StoreQueue.scala 103:23:@923.10]
  assign _T_2357 = offsetQ_8 < previousLoadHead; // @[StoreQueue.scala 103:75:@924.10]
  assign _T_2358 = _T_2356 & _T_2357; // @[StoreQueue.scala 103:49:@925.10]
  assign _T_2360 = _T_2358 == 1'h0; // @[StoreQueue.scala 103:9:@926.10]
  assign _T_2361 = _T_2115 & _T_2360; // @[StoreQueue.scala 102:49:@927.10]
  assign _GEN_720 = _T_2361 ? 1'h0 : checkBits_8; // @[StoreQueue.scala 103:96:@928.10]
  assign _GEN_721 = _T_2353 ? 1'h0 : _GEN_720; // @[StoreQueue.scala 100:102:@918.8]
  assign _GEN_722 = io_loadEmpty ? 1'h0 : _GEN_721; // @[StoreQueue.scala 98:26:@911.6]
  assign _GEN_723 = initBits_8 ? _T_2349 : _GEN_722; // @[StoreQueue.scala 94:35:@896.4]
  assign _T_2374 = _GEN_321 + 4'h1; // @[util.scala 10:8:@939.6]
  assign _GEN_424 = _T_2374 % 5'h10; // @[util.scala 10:14:@940.6]
  assign _T_2375 = _GEN_424[4:0]; // @[util.scala 10:14:@940.6]
  assign _T_2376 = _T_2375 == _GEN_1267; // @[StoreQueue.scala 96:56:@941.6]
  assign _T_2377 = io_loadEmpty & _T_2376; // @[StoreQueue.scala 95:50:@942.6]
  assign _T_2379 = _T_2377 == 1'h0; // @[StoreQueue.scala 95:35:@943.6]
  assign _T_2381 = previousLoadHead <= offsetQ_9; // @[StoreQueue.scala 100:35:@951.8]
  assign _T_2382 = offsetQ_9 < io_loadHead; // @[StoreQueue.scala 100:87:@952.8]
  assign _T_2383 = _T_2381 & _T_2382; // @[StoreQueue.scala 100:61:@953.8]
  assign _T_2386 = io_loadHead <= offsetQ_9; // @[StoreQueue.scala 103:23:@959.10]
  assign _T_2387 = offsetQ_9 < previousLoadHead; // @[StoreQueue.scala 103:75:@960.10]
  assign _T_2388 = _T_2386 & _T_2387; // @[StoreQueue.scala 103:49:@961.10]
  assign _T_2390 = _T_2388 == 1'h0; // @[StoreQueue.scala 103:9:@962.10]
  assign _T_2391 = _T_2115 & _T_2390; // @[StoreQueue.scala 102:49:@963.10]
  assign _GEN_740 = _T_2391 ? 1'h0 : checkBits_9; // @[StoreQueue.scala 103:96:@964.10]
  assign _GEN_741 = _T_2383 ? 1'h0 : _GEN_740; // @[StoreQueue.scala 100:102:@954.8]
  assign _GEN_742 = io_loadEmpty ? 1'h0 : _GEN_741; // @[StoreQueue.scala 98:26:@947.6]
  assign _GEN_743 = initBits_9 ? _T_2379 : _GEN_742; // @[StoreQueue.scala 94:35:@932.4]
  assign _T_2404 = _GEN_355 + 4'h1; // @[util.scala 10:8:@975.6]
  assign _GEN_442 = _T_2404 % 5'h10; // @[util.scala 10:14:@976.6]
  assign _T_2405 = _GEN_442[4:0]; // @[util.scala 10:14:@976.6]
  assign _T_2406 = _T_2405 == _GEN_1267; // @[StoreQueue.scala 96:56:@977.6]
  assign _T_2407 = io_loadEmpty & _T_2406; // @[StoreQueue.scala 95:50:@978.6]
  assign _T_2409 = _T_2407 == 1'h0; // @[StoreQueue.scala 95:35:@979.6]
  assign _T_2411 = previousLoadHead <= offsetQ_10; // @[StoreQueue.scala 100:35:@987.8]
  assign _T_2412 = offsetQ_10 < io_loadHead; // @[StoreQueue.scala 100:87:@988.8]
  assign _T_2413 = _T_2411 & _T_2412; // @[StoreQueue.scala 100:61:@989.8]
  assign _T_2416 = io_loadHead <= offsetQ_10; // @[StoreQueue.scala 103:23:@995.10]
  assign _T_2417 = offsetQ_10 < previousLoadHead; // @[StoreQueue.scala 103:75:@996.10]
  assign _T_2418 = _T_2416 & _T_2417; // @[StoreQueue.scala 103:49:@997.10]
  assign _T_2420 = _T_2418 == 1'h0; // @[StoreQueue.scala 103:9:@998.10]
  assign _T_2421 = _T_2115 & _T_2420; // @[StoreQueue.scala 102:49:@999.10]
  assign _GEN_760 = _T_2421 ? 1'h0 : checkBits_10; // @[StoreQueue.scala 103:96:@1000.10]
  assign _GEN_761 = _T_2413 ? 1'h0 : _GEN_760; // @[StoreQueue.scala 100:102:@990.8]
  assign _GEN_762 = io_loadEmpty ? 1'h0 : _GEN_761; // @[StoreQueue.scala 98:26:@983.6]
  assign _GEN_763 = initBits_10 ? _T_2409 : _GEN_762; // @[StoreQueue.scala 94:35:@968.4]
  assign _T_2434 = _GEN_389 + 4'h1; // @[util.scala 10:8:@1011.6]
  assign _GEN_458 = _T_2434 % 5'h10; // @[util.scala 10:14:@1012.6]
  assign _T_2435 = _GEN_458[4:0]; // @[util.scala 10:14:@1012.6]
  assign _T_2436 = _T_2435 == _GEN_1267; // @[StoreQueue.scala 96:56:@1013.6]
  assign _T_2437 = io_loadEmpty & _T_2436; // @[StoreQueue.scala 95:50:@1014.6]
  assign _T_2439 = _T_2437 == 1'h0; // @[StoreQueue.scala 95:35:@1015.6]
  assign _T_2441 = previousLoadHead <= offsetQ_11; // @[StoreQueue.scala 100:35:@1023.8]
  assign _T_2442 = offsetQ_11 < io_loadHead; // @[StoreQueue.scala 100:87:@1024.8]
  assign _T_2443 = _T_2441 & _T_2442; // @[StoreQueue.scala 100:61:@1025.8]
  assign _T_2446 = io_loadHead <= offsetQ_11; // @[StoreQueue.scala 103:23:@1031.10]
  assign _T_2447 = offsetQ_11 < previousLoadHead; // @[StoreQueue.scala 103:75:@1032.10]
  assign _T_2448 = _T_2446 & _T_2447; // @[StoreQueue.scala 103:49:@1033.10]
  assign _T_2450 = _T_2448 == 1'h0; // @[StoreQueue.scala 103:9:@1034.10]
  assign _T_2451 = _T_2115 & _T_2450; // @[StoreQueue.scala 102:49:@1035.10]
  assign _GEN_780 = _T_2451 ? 1'h0 : checkBits_11; // @[StoreQueue.scala 103:96:@1036.10]
  assign _GEN_781 = _T_2443 ? 1'h0 : _GEN_780; // @[StoreQueue.scala 100:102:@1026.8]
  assign _GEN_782 = io_loadEmpty ? 1'h0 : _GEN_781; // @[StoreQueue.scala 98:26:@1019.6]
  assign _GEN_783 = initBits_11 ? _T_2439 : _GEN_782; // @[StoreQueue.scala 94:35:@1004.4]
  assign _T_2464 = _GEN_423 + 4'h1; // @[util.scala 10:8:@1047.6]
  assign _GEN_476 = _T_2464 % 5'h10; // @[util.scala 10:14:@1048.6]
  assign _T_2465 = _GEN_476[4:0]; // @[util.scala 10:14:@1048.6]
  assign _T_2466 = _T_2465 == _GEN_1267; // @[StoreQueue.scala 96:56:@1049.6]
  assign _T_2467 = io_loadEmpty & _T_2466; // @[StoreQueue.scala 95:50:@1050.6]
  assign _T_2469 = _T_2467 == 1'h0; // @[StoreQueue.scala 95:35:@1051.6]
  assign _T_2471 = previousLoadHead <= offsetQ_12; // @[StoreQueue.scala 100:35:@1059.8]
  assign _T_2472 = offsetQ_12 < io_loadHead; // @[StoreQueue.scala 100:87:@1060.8]
  assign _T_2473 = _T_2471 & _T_2472; // @[StoreQueue.scala 100:61:@1061.8]
  assign _T_2476 = io_loadHead <= offsetQ_12; // @[StoreQueue.scala 103:23:@1067.10]
  assign _T_2477 = offsetQ_12 < previousLoadHead; // @[StoreQueue.scala 103:75:@1068.10]
  assign _T_2478 = _T_2476 & _T_2477; // @[StoreQueue.scala 103:49:@1069.10]
  assign _T_2480 = _T_2478 == 1'h0; // @[StoreQueue.scala 103:9:@1070.10]
  assign _T_2481 = _T_2115 & _T_2480; // @[StoreQueue.scala 102:49:@1071.10]
  assign _GEN_800 = _T_2481 ? 1'h0 : checkBits_12; // @[StoreQueue.scala 103:96:@1072.10]
  assign _GEN_801 = _T_2473 ? 1'h0 : _GEN_800; // @[StoreQueue.scala 100:102:@1062.8]
  assign _GEN_802 = io_loadEmpty ? 1'h0 : _GEN_801; // @[StoreQueue.scala 98:26:@1055.6]
  assign _GEN_803 = initBits_12 ? _T_2469 : _GEN_802; // @[StoreQueue.scala 94:35:@1040.4]
  assign _T_2494 = _GEN_457 + 4'h1; // @[util.scala 10:8:@1083.6]
  assign _GEN_492 = _T_2494 % 5'h10; // @[util.scala 10:14:@1084.6]
  assign _T_2495 = _GEN_492[4:0]; // @[util.scala 10:14:@1084.6]
  assign _T_2496 = _T_2495 == _GEN_1267; // @[StoreQueue.scala 96:56:@1085.6]
  assign _T_2497 = io_loadEmpty & _T_2496; // @[StoreQueue.scala 95:50:@1086.6]
  assign _T_2499 = _T_2497 == 1'h0; // @[StoreQueue.scala 95:35:@1087.6]
  assign _T_2501 = previousLoadHead <= offsetQ_13; // @[StoreQueue.scala 100:35:@1095.8]
  assign _T_2502 = offsetQ_13 < io_loadHead; // @[StoreQueue.scala 100:87:@1096.8]
  assign _T_2503 = _T_2501 & _T_2502; // @[StoreQueue.scala 100:61:@1097.8]
  assign _T_2506 = io_loadHead <= offsetQ_13; // @[StoreQueue.scala 103:23:@1103.10]
  assign _T_2507 = offsetQ_13 < previousLoadHead; // @[StoreQueue.scala 103:75:@1104.10]
  assign _T_2508 = _T_2506 & _T_2507; // @[StoreQueue.scala 103:49:@1105.10]
  assign _T_2510 = _T_2508 == 1'h0; // @[StoreQueue.scala 103:9:@1106.10]
  assign _T_2511 = _T_2115 & _T_2510; // @[StoreQueue.scala 102:49:@1107.10]
  assign _GEN_820 = _T_2511 ? 1'h0 : checkBits_13; // @[StoreQueue.scala 103:96:@1108.10]
  assign _GEN_821 = _T_2503 ? 1'h0 : _GEN_820; // @[StoreQueue.scala 100:102:@1098.8]
  assign _GEN_822 = io_loadEmpty ? 1'h0 : _GEN_821; // @[StoreQueue.scala 98:26:@1091.6]
  assign _GEN_823 = initBits_13 ? _T_2499 : _GEN_822; // @[StoreQueue.scala 94:35:@1076.4]
  assign _T_2524 = _GEN_491 + 4'h1; // @[util.scala 10:8:@1119.6]
  assign _GEN_510 = _T_2524 % 5'h10; // @[util.scala 10:14:@1120.6]
  assign _T_2525 = _GEN_510[4:0]; // @[util.scala 10:14:@1120.6]
  assign _T_2526 = _T_2525 == _GEN_1267; // @[StoreQueue.scala 96:56:@1121.6]
  assign _T_2527 = io_loadEmpty & _T_2526; // @[StoreQueue.scala 95:50:@1122.6]
  assign _T_2529 = _T_2527 == 1'h0; // @[StoreQueue.scala 95:35:@1123.6]
  assign _T_2531 = previousLoadHead <= offsetQ_14; // @[StoreQueue.scala 100:35:@1131.8]
  assign _T_2532 = offsetQ_14 < io_loadHead; // @[StoreQueue.scala 100:87:@1132.8]
  assign _T_2533 = _T_2531 & _T_2532; // @[StoreQueue.scala 100:61:@1133.8]
  assign _T_2536 = io_loadHead <= offsetQ_14; // @[StoreQueue.scala 103:23:@1139.10]
  assign _T_2537 = offsetQ_14 < previousLoadHead; // @[StoreQueue.scala 103:75:@1140.10]
  assign _T_2538 = _T_2536 & _T_2537; // @[StoreQueue.scala 103:49:@1141.10]
  assign _T_2540 = _T_2538 == 1'h0; // @[StoreQueue.scala 103:9:@1142.10]
  assign _T_2541 = _T_2115 & _T_2540; // @[StoreQueue.scala 102:49:@1143.10]
  assign _GEN_840 = _T_2541 ? 1'h0 : checkBits_14; // @[StoreQueue.scala 103:96:@1144.10]
  assign _GEN_841 = _T_2533 ? 1'h0 : _GEN_840; // @[StoreQueue.scala 100:102:@1134.8]
  assign _GEN_842 = io_loadEmpty ? 1'h0 : _GEN_841; // @[StoreQueue.scala 98:26:@1127.6]
  assign _GEN_843 = initBits_14 ? _T_2529 : _GEN_842; // @[StoreQueue.scala 94:35:@1112.4]
  assign _T_2554 = _GEN_525 + 4'h1; // @[util.scala 10:8:@1155.6]
  assign _GEN_526 = _T_2554 % 5'h10; // @[util.scala 10:14:@1156.6]
  assign _T_2555 = _GEN_526[4:0]; // @[util.scala 10:14:@1156.6]
  assign _T_2556 = _T_2555 == _GEN_1267; // @[StoreQueue.scala 96:56:@1157.6]
  assign _T_2557 = io_loadEmpty & _T_2556; // @[StoreQueue.scala 95:50:@1158.6]
  assign _T_2559 = _T_2557 == 1'h0; // @[StoreQueue.scala 95:35:@1159.6]
  assign _T_2561 = previousLoadHead <= offsetQ_15; // @[StoreQueue.scala 100:35:@1167.8]
  assign _T_2562 = offsetQ_15 < io_loadHead; // @[StoreQueue.scala 100:87:@1168.8]
  assign _T_2563 = _T_2561 & _T_2562; // @[StoreQueue.scala 100:61:@1169.8]
  assign _T_2566 = io_loadHead <= offsetQ_15; // @[StoreQueue.scala 103:23:@1175.10]
  assign _T_2567 = offsetQ_15 < previousLoadHead; // @[StoreQueue.scala 103:75:@1176.10]
  assign _T_2568 = _T_2566 & _T_2567; // @[StoreQueue.scala 103:49:@1177.10]
  assign _T_2570 = _T_2568 == 1'h0; // @[StoreQueue.scala 103:9:@1178.10]
  assign _T_2571 = _T_2115 & _T_2570; // @[StoreQueue.scala 102:49:@1179.10]
  assign _GEN_860 = _T_2571 ? 1'h0 : checkBits_15; // @[StoreQueue.scala 103:96:@1180.10]
  assign _GEN_861 = _T_2563 ? 1'h0 : _GEN_860; // @[StoreQueue.scala 100:102:@1170.8]
  assign _GEN_862 = io_loadEmpty ? 1'h0 : _GEN_861; // @[StoreQueue.scala 98:26:@1163.6]
  assign _GEN_863 = initBits_15 ? _T_2559 : _GEN_862; // @[StoreQueue.scala 94:35:@1148.4]
  assign _T_2573 = io_loadHead < io_loadTail; // @[StoreQueue.scala 119:103:@1184.4]
  assign _T_2575 = io_loadHead <= 4'h0; // @[StoreQueue.scala 120:17:@1185.4]
  assign _T_2577 = 4'h0 < io_loadTail; // @[StoreQueue.scala 120:35:@1186.4]
  assign _T_2578 = _T_2575 & _T_2577; // @[StoreQueue.scala 120:26:@1187.4]
  assign _T_2580 = io_loadEmpty == 1'h0; // @[StoreQueue.scala 120:50:@1188.4]
  assign _T_2582 = io_loadTail <= 4'h0; // @[StoreQueue.scala 120:81:@1189.4]
  assign _T_2584 = 4'h0 < io_loadHead; // @[StoreQueue.scala 120:99:@1190.4]
  assign _T_2585 = _T_2582 & _T_2584; // @[StoreQueue.scala 120:90:@1191.4]
  assign _T_2587 = _T_2585 == 1'h0; // @[StoreQueue.scala 120:67:@1192.4]
  assign _T_2588 = _T_2580 & _T_2587; // @[StoreQueue.scala 120:64:@1193.4]
  assign validEntriesInLoadQ_0 = _T_2573 ? _T_2578 : _T_2588; // @[StoreQueue.scala 119:90:@1194.4]
  assign _T_2592 = io_loadHead <= 4'h1; // @[StoreQueue.scala 120:17:@1196.4]
  assign _T_2594 = 4'h1 < io_loadTail; // @[StoreQueue.scala 120:35:@1197.4]
  assign _T_2595 = _T_2592 & _T_2594; // @[StoreQueue.scala 120:26:@1198.4]
  assign _T_2599 = io_loadTail <= 4'h1; // @[StoreQueue.scala 120:81:@1200.4]
  assign _T_2601 = 4'h1 < io_loadHead; // @[StoreQueue.scala 120:99:@1201.4]
  assign _T_2602 = _T_2599 & _T_2601; // @[StoreQueue.scala 120:90:@1202.4]
  assign _T_2604 = _T_2602 == 1'h0; // @[StoreQueue.scala 120:67:@1203.4]
  assign _T_2605 = _T_2580 & _T_2604; // @[StoreQueue.scala 120:64:@1204.4]
  assign validEntriesInLoadQ_1 = _T_2573 ? _T_2595 : _T_2605; // @[StoreQueue.scala 119:90:@1205.4]
  assign _T_2609 = io_loadHead <= 4'h2; // @[StoreQueue.scala 120:17:@1207.4]
  assign _T_2611 = 4'h2 < io_loadTail; // @[StoreQueue.scala 120:35:@1208.4]
  assign _T_2612 = _T_2609 & _T_2611; // @[StoreQueue.scala 120:26:@1209.4]
  assign _T_2616 = io_loadTail <= 4'h2; // @[StoreQueue.scala 120:81:@1211.4]
  assign _T_2618 = 4'h2 < io_loadHead; // @[StoreQueue.scala 120:99:@1212.4]
  assign _T_2619 = _T_2616 & _T_2618; // @[StoreQueue.scala 120:90:@1213.4]
  assign _T_2621 = _T_2619 == 1'h0; // @[StoreQueue.scala 120:67:@1214.4]
  assign _T_2622 = _T_2580 & _T_2621; // @[StoreQueue.scala 120:64:@1215.4]
  assign validEntriesInLoadQ_2 = _T_2573 ? _T_2612 : _T_2622; // @[StoreQueue.scala 119:90:@1216.4]
  assign _T_2626 = io_loadHead <= 4'h3; // @[StoreQueue.scala 120:17:@1218.4]
  assign _T_2628 = 4'h3 < io_loadTail; // @[StoreQueue.scala 120:35:@1219.4]
  assign _T_2629 = _T_2626 & _T_2628; // @[StoreQueue.scala 120:26:@1220.4]
  assign _T_2633 = io_loadTail <= 4'h3; // @[StoreQueue.scala 120:81:@1222.4]
  assign _T_2635 = 4'h3 < io_loadHead; // @[StoreQueue.scala 120:99:@1223.4]
  assign _T_2636 = _T_2633 & _T_2635; // @[StoreQueue.scala 120:90:@1224.4]
  assign _T_2638 = _T_2636 == 1'h0; // @[StoreQueue.scala 120:67:@1225.4]
  assign _T_2639 = _T_2580 & _T_2638; // @[StoreQueue.scala 120:64:@1226.4]
  assign validEntriesInLoadQ_3 = _T_2573 ? _T_2629 : _T_2639; // @[StoreQueue.scala 119:90:@1227.4]
  assign _T_2643 = io_loadHead <= 4'h4; // @[StoreQueue.scala 120:17:@1229.4]
  assign _T_2645 = 4'h4 < io_loadTail; // @[StoreQueue.scala 120:35:@1230.4]
  assign _T_2646 = _T_2643 & _T_2645; // @[StoreQueue.scala 120:26:@1231.4]
  assign _T_2650 = io_loadTail <= 4'h4; // @[StoreQueue.scala 120:81:@1233.4]
  assign _T_2652 = 4'h4 < io_loadHead; // @[StoreQueue.scala 120:99:@1234.4]
  assign _T_2653 = _T_2650 & _T_2652; // @[StoreQueue.scala 120:90:@1235.4]
  assign _T_2655 = _T_2653 == 1'h0; // @[StoreQueue.scala 120:67:@1236.4]
  assign _T_2656 = _T_2580 & _T_2655; // @[StoreQueue.scala 120:64:@1237.4]
  assign validEntriesInLoadQ_4 = _T_2573 ? _T_2646 : _T_2656; // @[StoreQueue.scala 119:90:@1238.4]
  assign _T_2660 = io_loadHead <= 4'h5; // @[StoreQueue.scala 120:17:@1240.4]
  assign _T_2662 = 4'h5 < io_loadTail; // @[StoreQueue.scala 120:35:@1241.4]
  assign _T_2663 = _T_2660 & _T_2662; // @[StoreQueue.scala 120:26:@1242.4]
  assign _T_2667 = io_loadTail <= 4'h5; // @[StoreQueue.scala 120:81:@1244.4]
  assign _T_2669 = 4'h5 < io_loadHead; // @[StoreQueue.scala 120:99:@1245.4]
  assign _T_2670 = _T_2667 & _T_2669; // @[StoreQueue.scala 120:90:@1246.4]
  assign _T_2672 = _T_2670 == 1'h0; // @[StoreQueue.scala 120:67:@1247.4]
  assign _T_2673 = _T_2580 & _T_2672; // @[StoreQueue.scala 120:64:@1248.4]
  assign validEntriesInLoadQ_5 = _T_2573 ? _T_2663 : _T_2673; // @[StoreQueue.scala 119:90:@1249.4]
  assign _T_2677 = io_loadHead <= 4'h6; // @[StoreQueue.scala 120:17:@1251.4]
  assign _T_2679 = 4'h6 < io_loadTail; // @[StoreQueue.scala 120:35:@1252.4]
  assign _T_2680 = _T_2677 & _T_2679; // @[StoreQueue.scala 120:26:@1253.4]
  assign _T_2684 = io_loadTail <= 4'h6; // @[StoreQueue.scala 120:81:@1255.4]
  assign _T_2686 = 4'h6 < io_loadHead; // @[StoreQueue.scala 120:99:@1256.4]
  assign _T_2687 = _T_2684 & _T_2686; // @[StoreQueue.scala 120:90:@1257.4]
  assign _T_2689 = _T_2687 == 1'h0; // @[StoreQueue.scala 120:67:@1258.4]
  assign _T_2690 = _T_2580 & _T_2689; // @[StoreQueue.scala 120:64:@1259.4]
  assign validEntriesInLoadQ_6 = _T_2573 ? _T_2680 : _T_2690; // @[StoreQueue.scala 119:90:@1260.4]
  assign _T_2694 = io_loadHead <= 4'h7; // @[StoreQueue.scala 120:17:@1262.4]
  assign _T_2696 = 4'h7 < io_loadTail; // @[StoreQueue.scala 120:35:@1263.4]
  assign _T_2697 = _T_2694 & _T_2696; // @[StoreQueue.scala 120:26:@1264.4]
  assign _T_2701 = io_loadTail <= 4'h7; // @[StoreQueue.scala 120:81:@1266.4]
  assign _T_2703 = 4'h7 < io_loadHead; // @[StoreQueue.scala 120:99:@1267.4]
  assign _T_2704 = _T_2701 & _T_2703; // @[StoreQueue.scala 120:90:@1268.4]
  assign _T_2706 = _T_2704 == 1'h0; // @[StoreQueue.scala 120:67:@1269.4]
  assign _T_2707 = _T_2580 & _T_2706; // @[StoreQueue.scala 120:64:@1270.4]
  assign validEntriesInLoadQ_7 = _T_2573 ? _T_2697 : _T_2707; // @[StoreQueue.scala 119:90:@1271.4]
  assign _T_2711 = io_loadHead <= 4'h8; // @[StoreQueue.scala 120:17:@1273.4]
  assign _T_2713 = 4'h8 < io_loadTail; // @[StoreQueue.scala 120:35:@1274.4]
  assign _T_2714 = _T_2711 & _T_2713; // @[StoreQueue.scala 120:26:@1275.4]
  assign _T_2718 = io_loadTail <= 4'h8; // @[StoreQueue.scala 120:81:@1277.4]
  assign _T_2720 = 4'h8 < io_loadHead; // @[StoreQueue.scala 120:99:@1278.4]
  assign _T_2721 = _T_2718 & _T_2720; // @[StoreQueue.scala 120:90:@1279.4]
  assign _T_2723 = _T_2721 == 1'h0; // @[StoreQueue.scala 120:67:@1280.4]
  assign _T_2724 = _T_2580 & _T_2723; // @[StoreQueue.scala 120:64:@1281.4]
  assign validEntriesInLoadQ_8 = _T_2573 ? _T_2714 : _T_2724; // @[StoreQueue.scala 119:90:@1282.4]
  assign _T_2728 = io_loadHead <= 4'h9; // @[StoreQueue.scala 120:17:@1284.4]
  assign _T_2730 = 4'h9 < io_loadTail; // @[StoreQueue.scala 120:35:@1285.4]
  assign _T_2731 = _T_2728 & _T_2730; // @[StoreQueue.scala 120:26:@1286.4]
  assign _T_2735 = io_loadTail <= 4'h9; // @[StoreQueue.scala 120:81:@1288.4]
  assign _T_2737 = 4'h9 < io_loadHead; // @[StoreQueue.scala 120:99:@1289.4]
  assign _T_2738 = _T_2735 & _T_2737; // @[StoreQueue.scala 120:90:@1290.4]
  assign _T_2740 = _T_2738 == 1'h0; // @[StoreQueue.scala 120:67:@1291.4]
  assign _T_2741 = _T_2580 & _T_2740; // @[StoreQueue.scala 120:64:@1292.4]
  assign validEntriesInLoadQ_9 = _T_2573 ? _T_2731 : _T_2741; // @[StoreQueue.scala 119:90:@1293.4]
  assign _T_2745 = io_loadHead <= 4'ha; // @[StoreQueue.scala 120:17:@1295.4]
  assign _T_2747 = 4'ha < io_loadTail; // @[StoreQueue.scala 120:35:@1296.4]
  assign _T_2748 = _T_2745 & _T_2747; // @[StoreQueue.scala 120:26:@1297.4]
  assign _T_2752 = io_loadTail <= 4'ha; // @[StoreQueue.scala 120:81:@1299.4]
  assign _T_2754 = 4'ha < io_loadHead; // @[StoreQueue.scala 120:99:@1300.4]
  assign _T_2755 = _T_2752 & _T_2754; // @[StoreQueue.scala 120:90:@1301.4]
  assign _T_2757 = _T_2755 == 1'h0; // @[StoreQueue.scala 120:67:@1302.4]
  assign _T_2758 = _T_2580 & _T_2757; // @[StoreQueue.scala 120:64:@1303.4]
  assign validEntriesInLoadQ_10 = _T_2573 ? _T_2748 : _T_2758; // @[StoreQueue.scala 119:90:@1304.4]
  assign _T_2762 = io_loadHead <= 4'hb; // @[StoreQueue.scala 120:17:@1306.4]
  assign _T_2764 = 4'hb < io_loadTail; // @[StoreQueue.scala 120:35:@1307.4]
  assign _T_2765 = _T_2762 & _T_2764; // @[StoreQueue.scala 120:26:@1308.4]
  assign _T_2769 = io_loadTail <= 4'hb; // @[StoreQueue.scala 120:81:@1310.4]
  assign _T_2771 = 4'hb < io_loadHead; // @[StoreQueue.scala 120:99:@1311.4]
  assign _T_2772 = _T_2769 & _T_2771; // @[StoreQueue.scala 120:90:@1312.4]
  assign _T_2774 = _T_2772 == 1'h0; // @[StoreQueue.scala 120:67:@1313.4]
  assign _T_2775 = _T_2580 & _T_2774; // @[StoreQueue.scala 120:64:@1314.4]
  assign validEntriesInLoadQ_11 = _T_2573 ? _T_2765 : _T_2775; // @[StoreQueue.scala 119:90:@1315.4]
  assign _T_2779 = io_loadHead <= 4'hc; // @[StoreQueue.scala 120:17:@1317.4]
  assign _T_2781 = 4'hc < io_loadTail; // @[StoreQueue.scala 120:35:@1318.4]
  assign _T_2782 = _T_2779 & _T_2781; // @[StoreQueue.scala 120:26:@1319.4]
  assign _T_2786 = io_loadTail <= 4'hc; // @[StoreQueue.scala 120:81:@1321.4]
  assign _T_2788 = 4'hc < io_loadHead; // @[StoreQueue.scala 120:99:@1322.4]
  assign _T_2789 = _T_2786 & _T_2788; // @[StoreQueue.scala 120:90:@1323.4]
  assign _T_2791 = _T_2789 == 1'h0; // @[StoreQueue.scala 120:67:@1324.4]
  assign _T_2792 = _T_2580 & _T_2791; // @[StoreQueue.scala 120:64:@1325.4]
  assign validEntriesInLoadQ_12 = _T_2573 ? _T_2782 : _T_2792; // @[StoreQueue.scala 119:90:@1326.4]
  assign _T_2796 = io_loadHead <= 4'hd; // @[StoreQueue.scala 120:17:@1328.4]
  assign _T_2798 = 4'hd < io_loadTail; // @[StoreQueue.scala 120:35:@1329.4]
  assign _T_2799 = _T_2796 & _T_2798; // @[StoreQueue.scala 120:26:@1330.4]
  assign _T_2803 = io_loadTail <= 4'hd; // @[StoreQueue.scala 120:81:@1332.4]
  assign _T_2805 = 4'hd < io_loadHead; // @[StoreQueue.scala 120:99:@1333.4]
  assign _T_2806 = _T_2803 & _T_2805; // @[StoreQueue.scala 120:90:@1334.4]
  assign _T_2808 = _T_2806 == 1'h0; // @[StoreQueue.scala 120:67:@1335.4]
  assign _T_2809 = _T_2580 & _T_2808; // @[StoreQueue.scala 120:64:@1336.4]
  assign validEntriesInLoadQ_13 = _T_2573 ? _T_2799 : _T_2809; // @[StoreQueue.scala 119:90:@1337.4]
  assign _T_2813 = io_loadHead <= 4'he; // @[StoreQueue.scala 120:17:@1339.4]
  assign _T_2815 = 4'he < io_loadTail; // @[StoreQueue.scala 120:35:@1340.4]
  assign _T_2816 = _T_2813 & _T_2815; // @[StoreQueue.scala 120:26:@1341.4]
  assign _T_2820 = io_loadTail <= 4'he; // @[StoreQueue.scala 120:81:@1343.4]
  assign _T_2822 = 4'he < io_loadHead; // @[StoreQueue.scala 120:99:@1344.4]
  assign _T_2823 = _T_2820 & _T_2822; // @[StoreQueue.scala 120:90:@1345.4]
  assign _T_2825 = _T_2823 == 1'h0; // @[StoreQueue.scala 120:67:@1346.4]
  assign _T_2826 = _T_2580 & _T_2825; // @[StoreQueue.scala 120:64:@1347.4]
  assign validEntriesInLoadQ_14 = _T_2573 ? _T_2816 : _T_2826; // @[StoreQueue.scala 119:90:@1348.4]
  assign validEntriesInLoadQ_15 = _T_2573 ? 1'h0 : _T_2580; // @[StoreQueue.scala 119:90:@1359.4]
  assign _GEN_865 = 4'h1 == head ? offsetQ_1 : offsetQ_0; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_866 = 4'h2 == head ? offsetQ_2 : _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_867 = 4'h3 == head ? offsetQ_3 : _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_868 = 4'h4 == head ? offsetQ_4 : _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_869 = 4'h5 == head ? offsetQ_5 : _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_870 = 4'h6 == head ? offsetQ_6 : _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_871 = 4'h7 == head ? offsetQ_7 : _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_872 = 4'h8 == head ? offsetQ_8 : _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_873 = 4'h9 == head ? offsetQ_9 : _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_874 = 4'ha == head ? offsetQ_10 : _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_875 = 4'hb == head ? offsetQ_11 : _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_876 = 4'hc == head ? offsetQ_12 : _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_877 = 4'hd == head ? offsetQ_13 : _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_878 = 4'he == head ? offsetQ_14 : _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_879 = 4'hf == head ? offsetQ_15 : _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  assign _T_2869 = io_loadHead <= _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  assign loadsToCheck_0 = _T_2869 ? _T_2575 : 1'h1; // @[StoreQueue.scala 126:83:@1385.4]
  assign _T_2899 = 4'h1 <= _GEN_879; // @[StoreQueue.scala 127:37:@1388.4]
  assign _T_2900 = _T_2592 & _T_2899; // @[StoreQueue.scala 127:28:@1389.4]
  assign _T_2905 = _GEN_879 < 4'h1; // @[StoreQueue.scala 127:71:@1390.4]
  assign _T_2908 = _T_2905 & _T_2601; // @[StoreQueue.scala 127:79:@1392.4]
  assign _T_2910 = _T_2908 == 1'h0; // @[StoreQueue.scala 127:55:@1393.4]
  assign loadsToCheck_1 = _T_2869 ? _T_2900 : _T_2910; // @[StoreQueue.scala 126:83:@1394.4]
  assign _T_2922 = 4'h2 <= _GEN_879; // @[StoreQueue.scala 127:37:@1397.4]
  assign _T_2923 = _T_2609 & _T_2922; // @[StoreQueue.scala 127:28:@1398.4]
  assign _T_2928 = _GEN_879 < 4'h2; // @[StoreQueue.scala 127:71:@1399.4]
  assign _T_2931 = _T_2928 & _T_2618; // @[StoreQueue.scala 127:79:@1401.4]
  assign _T_2933 = _T_2931 == 1'h0; // @[StoreQueue.scala 127:55:@1402.4]
  assign loadsToCheck_2 = _T_2869 ? _T_2923 : _T_2933; // @[StoreQueue.scala 126:83:@1403.4]
  assign _T_2945 = 4'h3 <= _GEN_879; // @[StoreQueue.scala 127:37:@1406.4]
  assign _T_2946 = _T_2626 & _T_2945; // @[StoreQueue.scala 127:28:@1407.4]
  assign _T_2951 = _GEN_879 < 4'h3; // @[StoreQueue.scala 127:71:@1408.4]
  assign _T_2954 = _T_2951 & _T_2635; // @[StoreQueue.scala 127:79:@1410.4]
  assign _T_2956 = _T_2954 == 1'h0; // @[StoreQueue.scala 127:55:@1411.4]
  assign loadsToCheck_3 = _T_2869 ? _T_2946 : _T_2956; // @[StoreQueue.scala 126:83:@1412.4]
  assign _T_2968 = 4'h4 <= _GEN_879; // @[StoreQueue.scala 127:37:@1415.4]
  assign _T_2969 = _T_2643 & _T_2968; // @[StoreQueue.scala 127:28:@1416.4]
  assign _T_2974 = _GEN_879 < 4'h4; // @[StoreQueue.scala 127:71:@1417.4]
  assign _T_2977 = _T_2974 & _T_2652; // @[StoreQueue.scala 127:79:@1419.4]
  assign _T_2979 = _T_2977 == 1'h0; // @[StoreQueue.scala 127:55:@1420.4]
  assign loadsToCheck_4 = _T_2869 ? _T_2969 : _T_2979; // @[StoreQueue.scala 126:83:@1421.4]
  assign _T_2991 = 4'h5 <= _GEN_879; // @[StoreQueue.scala 127:37:@1424.4]
  assign _T_2992 = _T_2660 & _T_2991; // @[StoreQueue.scala 127:28:@1425.4]
  assign _T_2997 = _GEN_879 < 4'h5; // @[StoreQueue.scala 127:71:@1426.4]
  assign _T_3000 = _T_2997 & _T_2669; // @[StoreQueue.scala 127:79:@1428.4]
  assign _T_3002 = _T_3000 == 1'h0; // @[StoreQueue.scala 127:55:@1429.4]
  assign loadsToCheck_5 = _T_2869 ? _T_2992 : _T_3002; // @[StoreQueue.scala 126:83:@1430.4]
  assign _T_3014 = 4'h6 <= _GEN_879; // @[StoreQueue.scala 127:37:@1433.4]
  assign _T_3015 = _T_2677 & _T_3014; // @[StoreQueue.scala 127:28:@1434.4]
  assign _T_3020 = _GEN_879 < 4'h6; // @[StoreQueue.scala 127:71:@1435.4]
  assign _T_3023 = _T_3020 & _T_2686; // @[StoreQueue.scala 127:79:@1437.4]
  assign _T_3025 = _T_3023 == 1'h0; // @[StoreQueue.scala 127:55:@1438.4]
  assign loadsToCheck_6 = _T_2869 ? _T_3015 : _T_3025; // @[StoreQueue.scala 126:83:@1439.4]
  assign _T_3037 = 4'h7 <= _GEN_879; // @[StoreQueue.scala 127:37:@1442.4]
  assign _T_3038 = _T_2694 & _T_3037; // @[StoreQueue.scala 127:28:@1443.4]
  assign _T_3043 = _GEN_879 < 4'h7; // @[StoreQueue.scala 127:71:@1444.4]
  assign _T_3046 = _T_3043 & _T_2703; // @[StoreQueue.scala 127:79:@1446.4]
  assign _T_3048 = _T_3046 == 1'h0; // @[StoreQueue.scala 127:55:@1447.4]
  assign loadsToCheck_7 = _T_2869 ? _T_3038 : _T_3048; // @[StoreQueue.scala 126:83:@1448.4]
  assign _T_3060 = 4'h8 <= _GEN_879; // @[StoreQueue.scala 127:37:@1451.4]
  assign _T_3061 = _T_2711 & _T_3060; // @[StoreQueue.scala 127:28:@1452.4]
  assign _T_3066 = _GEN_879 < 4'h8; // @[StoreQueue.scala 127:71:@1453.4]
  assign _T_3069 = _T_3066 & _T_2720; // @[StoreQueue.scala 127:79:@1455.4]
  assign _T_3071 = _T_3069 == 1'h0; // @[StoreQueue.scala 127:55:@1456.4]
  assign loadsToCheck_8 = _T_2869 ? _T_3061 : _T_3071; // @[StoreQueue.scala 126:83:@1457.4]
  assign _T_3083 = 4'h9 <= _GEN_879; // @[StoreQueue.scala 127:37:@1460.4]
  assign _T_3084 = _T_2728 & _T_3083; // @[StoreQueue.scala 127:28:@1461.4]
  assign _T_3089 = _GEN_879 < 4'h9; // @[StoreQueue.scala 127:71:@1462.4]
  assign _T_3092 = _T_3089 & _T_2737; // @[StoreQueue.scala 127:79:@1464.4]
  assign _T_3094 = _T_3092 == 1'h0; // @[StoreQueue.scala 127:55:@1465.4]
  assign loadsToCheck_9 = _T_2869 ? _T_3084 : _T_3094; // @[StoreQueue.scala 126:83:@1466.4]
  assign _T_3106 = 4'ha <= _GEN_879; // @[StoreQueue.scala 127:37:@1469.4]
  assign _T_3107 = _T_2745 & _T_3106; // @[StoreQueue.scala 127:28:@1470.4]
  assign _T_3112 = _GEN_879 < 4'ha; // @[StoreQueue.scala 127:71:@1471.4]
  assign _T_3115 = _T_3112 & _T_2754; // @[StoreQueue.scala 127:79:@1473.4]
  assign _T_3117 = _T_3115 == 1'h0; // @[StoreQueue.scala 127:55:@1474.4]
  assign loadsToCheck_10 = _T_2869 ? _T_3107 : _T_3117; // @[StoreQueue.scala 126:83:@1475.4]
  assign _T_3129 = 4'hb <= _GEN_879; // @[StoreQueue.scala 127:37:@1478.4]
  assign _T_3130 = _T_2762 & _T_3129; // @[StoreQueue.scala 127:28:@1479.4]
  assign _T_3135 = _GEN_879 < 4'hb; // @[StoreQueue.scala 127:71:@1480.4]
  assign _T_3138 = _T_3135 & _T_2771; // @[StoreQueue.scala 127:79:@1482.4]
  assign _T_3140 = _T_3138 == 1'h0; // @[StoreQueue.scala 127:55:@1483.4]
  assign loadsToCheck_11 = _T_2869 ? _T_3130 : _T_3140; // @[StoreQueue.scala 126:83:@1484.4]
  assign _T_3152 = 4'hc <= _GEN_879; // @[StoreQueue.scala 127:37:@1487.4]
  assign _T_3153 = _T_2779 & _T_3152; // @[StoreQueue.scala 127:28:@1488.4]
  assign _T_3158 = _GEN_879 < 4'hc; // @[StoreQueue.scala 127:71:@1489.4]
  assign _T_3161 = _T_3158 & _T_2788; // @[StoreQueue.scala 127:79:@1491.4]
  assign _T_3163 = _T_3161 == 1'h0; // @[StoreQueue.scala 127:55:@1492.4]
  assign loadsToCheck_12 = _T_2869 ? _T_3153 : _T_3163; // @[StoreQueue.scala 126:83:@1493.4]
  assign _T_3175 = 4'hd <= _GEN_879; // @[StoreQueue.scala 127:37:@1496.4]
  assign _T_3176 = _T_2796 & _T_3175; // @[StoreQueue.scala 127:28:@1497.4]
  assign _T_3181 = _GEN_879 < 4'hd; // @[StoreQueue.scala 127:71:@1498.4]
  assign _T_3184 = _T_3181 & _T_2805; // @[StoreQueue.scala 127:79:@1500.4]
  assign _T_3186 = _T_3184 == 1'h0; // @[StoreQueue.scala 127:55:@1501.4]
  assign loadsToCheck_13 = _T_2869 ? _T_3176 : _T_3186; // @[StoreQueue.scala 126:83:@1502.4]
  assign _T_3198 = 4'he <= _GEN_879; // @[StoreQueue.scala 127:37:@1505.4]
  assign _T_3199 = _T_2813 & _T_3198; // @[StoreQueue.scala 127:28:@1506.4]
  assign _T_3204 = _GEN_879 < 4'he; // @[StoreQueue.scala 127:71:@1507.4]
  assign _T_3207 = _T_3204 & _T_2822; // @[StoreQueue.scala 127:79:@1509.4]
  assign _T_3209 = _T_3207 == 1'h0; // @[StoreQueue.scala 127:55:@1510.4]
  assign loadsToCheck_14 = _T_2869 ? _T_3199 : _T_3209; // @[StoreQueue.scala 126:83:@1511.4]
  assign _T_3221 = 4'hf <= _GEN_879; // @[StoreQueue.scala 127:37:@1514.4]
  assign loadsToCheck_15 = _T_2869 ? _T_3221 : 1'h1; // @[StoreQueue.scala 126:83:@1520.4]
  assign _T_3255 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[StoreQueue.scala 133:16:@1538.4]
  assign _GEN_881 = 4'h1 == head ? checkBits_1 : checkBits_0; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_882 = 4'h2 == head ? checkBits_2 : _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_883 = 4'h3 == head ? checkBits_3 : _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_884 = 4'h4 == head ? checkBits_4 : _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_885 = 4'h5 == head ? checkBits_5 : _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_886 = 4'h6 == head ? checkBits_6 : _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_887 = 4'h7 == head ? checkBits_7 : _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_888 = 4'h8 == head ? checkBits_8 : _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_889 = 4'h9 == head ? checkBits_9 : _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_890 = 4'ha == head ? checkBits_10 : _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_891 = 4'hb == head ? checkBits_11 : _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_892 = 4'hc == head ? checkBits_12 : _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_893 = 4'hd == head ? checkBits_13 : _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_894 = 4'he == head ? checkBits_14 : _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_895 = 4'hf == head ? checkBits_15 : _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  assign entriesToCheck_0 = _T_3255 & _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  assign _T_3260 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[StoreQueue.scala 133:16:@1540.4]
  assign entriesToCheck_1 = _T_3260 & _GEN_895; // @[StoreQueue.scala 133:24:@1541.4]
  assign _T_3265 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[StoreQueue.scala 133:16:@1542.4]
  assign entriesToCheck_2 = _T_3265 & _GEN_895; // @[StoreQueue.scala 133:24:@1543.4]
  assign _T_3270 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[StoreQueue.scala 133:16:@1544.4]
  assign entriesToCheck_3 = _T_3270 & _GEN_895; // @[StoreQueue.scala 133:24:@1545.4]
  assign _T_3275 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[StoreQueue.scala 133:16:@1546.4]
  assign entriesToCheck_4 = _T_3275 & _GEN_895; // @[StoreQueue.scala 133:24:@1547.4]
  assign _T_3280 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[StoreQueue.scala 133:16:@1548.4]
  assign entriesToCheck_5 = _T_3280 & _GEN_895; // @[StoreQueue.scala 133:24:@1549.4]
  assign _T_3285 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[StoreQueue.scala 133:16:@1550.4]
  assign entriesToCheck_6 = _T_3285 & _GEN_895; // @[StoreQueue.scala 133:24:@1551.4]
  assign _T_3290 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[StoreQueue.scala 133:16:@1552.4]
  assign entriesToCheck_7 = _T_3290 & _GEN_895; // @[StoreQueue.scala 133:24:@1553.4]
  assign _T_3295 = loadsToCheck_8 & validEntriesInLoadQ_8; // @[StoreQueue.scala 133:16:@1554.4]
  assign entriesToCheck_8 = _T_3295 & _GEN_895; // @[StoreQueue.scala 133:24:@1555.4]
  assign _T_3300 = loadsToCheck_9 & validEntriesInLoadQ_9; // @[StoreQueue.scala 133:16:@1556.4]
  assign entriesToCheck_9 = _T_3300 & _GEN_895; // @[StoreQueue.scala 133:24:@1557.4]
  assign _T_3305 = loadsToCheck_10 & validEntriesInLoadQ_10; // @[StoreQueue.scala 133:16:@1558.4]
  assign entriesToCheck_10 = _T_3305 & _GEN_895; // @[StoreQueue.scala 133:24:@1559.4]
  assign _T_3310 = loadsToCheck_11 & validEntriesInLoadQ_11; // @[StoreQueue.scala 133:16:@1560.4]
  assign entriesToCheck_11 = _T_3310 & _GEN_895; // @[StoreQueue.scala 133:24:@1561.4]
  assign _T_3315 = loadsToCheck_12 & validEntriesInLoadQ_12; // @[StoreQueue.scala 133:16:@1562.4]
  assign entriesToCheck_12 = _T_3315 & _GEN_895; // @[StoreQueue.scala 133:24:@1563.4]
  assign _T_3320 = loadsToCheck_13 & validEntriesInLoadQ_13; // @[StoreQueue.scala 133:16:@1564.4]
  assign entriesToCheck_13 = _T_3320 & _GEN_895; // @[StoreQueue.scala 133:24:@1565.4]
  assign _T_3325 = loadsToCheck_14 & validEntriesInLoadQ_14; // @[StoreQueue.scala 133:16:@1566.4]
  assign entriesToCheck_14 = _T_3325 & _GEN_895; // @[StoreQueue.scala 133:24:@1567.4]
  assign _T_3330 = loadsToCheck_15 & validEntriesInLoadQ_15; // @[StoreQueue.scala 133:16:@1568.4]
  assign entriesToCheck_15 = _T_3330 & _GEN_895; // @[StoreQueue.scala 133:24:@1569.4]
  assign _T_3378 = entriesToCheck_0 == 1'h0; // @[StoreQueue.scala 140:34:@1588.4]
  assign _T_3379 = _T_3378 | io_loadDataDone_0; // @[StoreQueue.scala 140:64:@1589.4]
  assign _GEN_897 = 4'h1 == head ? addrQ_1 : addrQ_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_898 = 4'h2 == head ? addrQ_2 : _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_899 = 4'h3 == head ? addrQ_3 : _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_900 = 4'h4 == head ? addrQ_4 : _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_901 = 4'h5 == head ? addrQ_5 : _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_902 = 4'h6 == head ? addrQ_6 : _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_903 = 4'h7 == head ? addrQ_7 : _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_904 = 4'h8 == head ? addrQ_8 : _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_905 = 4'h9 == head ? addrQ_9 : _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_906 = 4'ha == head ? addrQ_10 : _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_907 = 4'hb == head ? addrQ_11 : _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_908 = 4'hc == head ? addrQ_12 : _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_909 = 4'hd == head ? addrQ_13 : _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_910 = 4'he == head ? addrQ_14 : _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_911 = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3383 = _GEN_911 != io_loadAddressQueue_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3384 = io_loadAddressDone_0 & _T_3383; // @[StoreQueue.scala 141:36:@1591.4]
  assign noConflicts_0 = _T_3379 | _T_3384; // @[StoreQueue.scala 140:95:@1592.4]
  assign _T_3387 = entriesToCheck_1 == 1'h0; // @[StoreQueue.scala 140:34:@1594.4]
  assign _T_3388 = _T_3387 | io_loadDataDone_1; // @[StoreQueue.scala 140:64:@1595.4]
  assign _T_3392 = _GEN_911 != io_loadAddressQueue_1; // @[StoreQueue.scala 141:51:@1596.4]
  assign _T_3393 = io_loadAddressDone_1 & _T_3392; // @[StoreQueue.scala 141:36:@1597.4]
  assign noConflicts_1 = _T_3388 | _T_3393; // @[StoreQueue.scala 140:95:@1598.4]
  assign _T_3396 = entriesToCheck_2 == 1'h0; // @[StoreQueue.scala 140:34:@1600.4]
  assign _T_3397 = _T_3396 | io_loadDataDone_2; // @[StoreQueue.scala 140:64:@1601.4]
  assign _T_3401 = _GEN_911 != io_loadAddressQueue_2; // @[StoreQueue.scala 141:51:@1602.4]
  assign _T_3402 = io_loadAddressDone_2 & _T_3401; // @[StoreQueue.scala 141:36:@1603.4]
  assign noConflicts_2 = _T_3397 | _T_3402; // @[StoreQueue.scala 140:95:@1604.4]
  assign _T_3405 = entriesToCheck_3 == 1'h0; // @[StoreQueue.scala 140:34:@1606.4]
  assign _T_3406 = _T_3405 | io_loadDataDone_3; // @[StoreQueue.scala 140:64:@1607.4]
  assign _T_3410 = _GEN_911 != io_loadAddressQueue_3; // @[StoreQueue.scala 141:51:@1608.4]
  assign _T_3411 = io_loadAddressDone_3 & _T_3410; // @[StoreQueue.scala 141:36:@1609.4]
  assign noConflicts_3 = _T_3406 | _T_3411; // @[StoreQueue.scala 140:95:@1610.4]
  assign _T_3414 = entriesToCheck_4 == 1'h0; // @[StoreQueue.scala 140:34:@1612.4]
  assign _T_3415 = _T_3414 | io_loadDataDone_4; // @[StoreQueue.scala 140:64:@1613.4]
  assign _T_3419 = _GEN_911 != io_loadAddressQueue_4; // @[StoreQueue.scala 141:51:@1614.4]
  assign _T_3420 = io_loadAddressDone_4 & _T_3419; // @[StoreQueue.scala 141:36:@1615.4]
  assign noConflicts_4 = _T_3415 | _T_3420; // @[StoreQueue.scala 140:95:@1616.4]
  assign _T_3423 = entriesToCheck_5 == 1'h0; // @[StoreQueue.scala 140:34:@1618.4]
  assign _T_3424 = _T_3423 | io_loadDataDone_5; // @[StoreQueue.scala 140:64:@1619.4]
  assign _T_3428 = _GEN_911 != io_loadAddressQueue_5; // @[StoreQueue.scala 141:51:@1620.4]
  assign _T_3429 = io_loadAddressDone_5 & _T_3428; // @[StoreQueue.scala 141:36:@1621.4]
  assign noConflicts_5 = _T_3424 | _T_3429; // @[StoreQueue.scala 140:95:@1622.4]
  assign _T_3432 = entriesToCheck_6 == 1'h0; // @[StoreQueue.scala 140:34:@1624.4]
  assign _T_3433 = _T_3432 | io_loadDataDone_6; // @[StoreQueue.scala 140:64:@1625.4]
  assign _T_3437 = _GEN_911 != io_loadAddressQueue_6; // @[StoreQueue.scala 141:51:@1626.4]
  assign _T_3438 = io_loadAddressDone_6 & _T_3437; // @[StoreQueue.scala 141:36:@1627.4]
  assign noConflicts_6 = _T_3433 | _T_3438; // @[StoreQueue.scala 140:95:@1628.4]
  assign _T_3441 = entriesToCheck_7 == 1'h0; // @[StoreQueue.scala 140:34:@1630.4]
  assign _T_3442 = _T_3441 | io_loadDataDone_7; // @[StoreQueue.scala 140:64:@1631.4]
  assign _T_3446 = _GEN_911 != io_loadAddressQueue_7; // @[StoreQueue.scala 141:51:@1632.4]
  assign _T_3447 = io_loadAddressDone_7 & _T_3446; // @[StoreQueue.scala 141:36:@1633.4]
  assign noConflicts_7 = _T_3442 | _T_3447; // @[StoreQueue.scala 140:95:@1634.4]
  assign _T_3450 = entriesToCheck_8 == 1'h0; // @[StoreQueue.scala 140:34:@1636.4]
  assign _T_3451 = _T_3450 | io_loadDataDone_8; // @[StoreQueue.scala 140:64:@1637.4]
  assign _T_3455 = _GEN_911 != io_loadAddressQueue_8; // @[StoreQueue.scala 141:51:@1638.4]
  assign _T_3456 = io_loadAddressDone_8 & _T_3455; // @[StoreQueue.scala 141:36:@1639.4]
  assign noConflicts_8 = _T_3451 | _T_3456; // @[StoreQueue.scala 140:95:@1640.4]
  assign _T_3459 = entriesToCheck_9 == 1'h0; // @[StoreQueue.scala 140:34:@1642.4]
  assign _T_3460 = _T_3459 | io_loadDataDone_9; // @[StoreQueue.scala 140:64:@1643.4]
  assign _T_3464 = _GEN_911 != io_loadAddressQueue_9; // @[StoreQueue.scala 141:51:@1644.4]
  assign _T_3465 = io_loadAddressDone_9 & _T_3464; // @[StoreQueue.scala 141:36:@1645.4]
  assign noConflicts_9 = _T_3460 | _T_3465; // @[StoreQueue.scala 140:95:@1646.4]
  assign _T_3468 = entriesToCheck_10 == 1'h0; // @[StoreQueue.scala 140:34:@1648.4]
  assign _T_3469 = _T_3468 | io_loadDataDone_10; // @[StoreQueue.scala 140:64:@1649.4]
  assign _T_3473 = _GEN_911 != io_loadAddressQueue_10; // @[StoreQueue.scala 141:51:@1650.4]
  assign _T_3474 = io_loadAddressDone_10 & _T_3473; // @[StoreQueue.scala 141:36:@1651.4]
  assign noConflicts_10 = _T_3469 | _T_3474; // @[StoreQueue.scala 140:95:@1652.4]
  assign _T_3477 = entriesToCheck_11 == 1'h0; // @[StoreQueue.scala 140:34:@1654.4]
  assign _T_3478 = _T_3477 | io_loadDataDone_11; // @[StoreQueue.scala 140:64:@1655.4]
  assign _T_3482 = _GEN_911 != io_loadAddressQueue_11; // @[StoreQueue.scala 141:51:@1656.4]
  assign _T_3483 = io_loadAddressDone_11 & _T_3482; // @[StoreQueue.scala 141:36:@1657.4]
  assign noConflicts_11 = _T_3478 | _T_3483; // @[StoreQueue.scala 140:95:@1658.4]
  assign _T_3486 = entriesToCheck_12 == 1'h0; // @[StoreQueue.scala 140:34:@1660.4]
  assign _T_3487 = _T_3486 | io_loadDataDone_12; // @[StoreQueue.scala 140:64:@1661.4]
  assign _T_3491 = _GEN_911 != io_loadAddressQueue_12; // @[StoreQueue.scala 141:51:@1662.4]
  assign _T_3492 = io_loadAddressDone_12 & _T_3491; // @[StoreQueue.scala 141:36:@1663.4]
  assign noConflicts_12 = _T_3487 | _T_3492; // @[StoreQueue.scala 140:95:@1664.4]
  assign _T_3495 = entriesToCheck_13 == 1'h0; // @[StoreQueue.scala 140:34:@1666.4]
  assign _T_3496 = _T_3495 | io_loadDataDone_13; // @[StoreQueue.scala 140:64:@1667.4]
  assign _T_3500 = _GEN_911 != io_loadAddressQueue_13; // @[StoreQueue.scala 141:51:@1668.4]
  assign _T_3501 = io_loadAddressDone_13 & _T_3500; // @[StoreQueue.scala 141:36:@1669.4]
  assign noConflicts_13 = _T_3496 | _T_3501; // @[StoreQueue.scala 140:95:@1670.4]
  assign _T_3504 = entriesToCheck_14 == 1'h0; // @[StoreQueue.scala 140:34:@1672.4]
  assign _T_3505 = _T_3504 | io_loadDataDone_14; // @[StoreQueue.scala 140:64:@1673.4]
  assign _T_3509 = _GEN_911 != io_loadAddressQueue_14; // @[StoreQueue.scala 141:51:@1674.4]
  assign _T_3510 = io_loadAddressDone_14 & _T_3509; // @[StoreQueue.scala 141:36:@1675.4]
  assign noConflicts_14 = _T_3505 | _T_3510; // @[StoreQueue.scala 140:95:@1676.4]
  assign _T_3513 = entriesToCheck_15 == 1'h0; // @[StoreQueue.scala 140:34:@1678.4]
  assign _T_3514 = _T_3513 | io_loadDataDone_15; // @[StoreQueue.scala 140:64:@1679.4]
  assign _T_3518 = _GEN_911 != io_loadAddressQueue_15; // @[StoreQueue.scala 141:51:@1680.4]
  assign _T_3519 = io_loadAddressDone_15 & _T_3518; // @[StoreQueue.scala 141:36:@1681.4]
  assign noConflicts_15 = _T_3514 | _T_3519; // @[StoreQueue.scala 140:95:@1682.4]
  assign _GEN_913 = 4'h1 == head ? addrKnown_1 : addrKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_914 = 4'h2 == head ? addrKnown_2 : _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_915 = 4'h3 == head ? addrKnown_3 : _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_916 = 4'h4 == head ? addrKnown_4 : _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_917 = 4'h5 == head ? addrKnown_5 : _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_918 = 4'h6 == head ? addrKnown_6 : _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_919 = 4'h7 == head ? addrKnown_7 : _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_920 = 4'h8 == head ? addrKnown_8 : _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_921 = 4'h9 == head ? addrKnown_9 : _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_922 = 4'ha == head ? addrKnown_10 : _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_923 = 4'hb == head ? addrKnown_11 : _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_924 = 4'hc == head ? addrKnown_12 : _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_925 = 4'hd == head ? addrKnown_13 : _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_926 = 4'he == head ? addrKnown_14 : _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_927 = 4'hf == head ? addrKnown_15 : _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_929 = 4'h1 == head ? dataKnown_1 : dataKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_930 = 4'h2 == head ? dataKnown_2 : _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_931 = 4'h3 == head ? dataKnown_3 : _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_932 = 4'h4 == head ? dataKnown_4 : _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_933 = 4'h5 == head ? dataKnown_5 : _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_934 = 4'h6 == head ? dataKnown_6 : _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_935 = 4'h7 == head ? dataKnown_7 : _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_936 = 4'h8 == head ? dataKnown_8 : _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_937 = 4'h9 == head ? dataKnown_9 : _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_938 = 4'ha == head ? dataKnown_10 : _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_939 = 4'hb == head ? dataKnown_11 : _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_940 = 4'hc == head ? dataKnown_12 : _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_941 = 4'hd == head ? dataKnown_13 : _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_942 = 4'he == head ? dataKnown_14 : _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_943 = 4'hf == head ? dataKnown_15 : _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  assign _T_3527 = _GEN_927 & _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_945 = 4'h1 == head ? storeCompleted_1 : storeCompleted_0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_946 = 4'h2 == head ? storeCompleted_2 : _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_947 = 4'h3 == head ? storeCompleted_3 : _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_948 = 4'h4 == head ? storeCompleted_4 : _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_949 = 4'h5 == head ? storeCompleted_5 : _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_950 = 4'h6 == head ? storeCompleted_6 : _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_951 = 4'h7 == head ? storeCompleted_7 : _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_952 = 4'h8 == head ? storeCompleted_8 : _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_953 = 4'h9 == head ? storeCompleted_9 : _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_954 = 4'ha == head ? storeCompleted_10 : _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_955 = 4'hb == head ? storeCompleted_11 : _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_956 = 4'hc == head ? storeCompleted_12 : _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_957 = 4'hd == head ? storeCompleted_13 : _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_958 = 4'he == head ? storeCompleted_14 : _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_959 = 4'hf == head ? storeCompleted_15 : _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3532 = _GEN_959 == 1'h0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3533 = _T_3527 & _T_3532; // @[StoreQueue.scala 154:63:@1686.4]
  assign _T_3536 = noConflicts_0 & noConflicts_1; // @[StoreQueue.scala 154:109:@1688.4]
  assign _T_3537 = _T_3536 & noConflicts_2; // @[StoreQueue.scala 154:109:@1689.4]
  assign _T_3538 = _T_3537 & noConflicts_3; // @[StoreQueue.scala 154:109:@1690.4]
  assign _T_3539 = _T_3538 & noConflicts_4; // @[StoreQueue.scala 154:109:@1691.4]
  assign _T_3540 = _T_3539 & noConflicts_5; // @[StoreQueue.scala 154:109:@1692.4]
  assign _T_3541 = _T_3540 & noConflicts_6; // @[StoreQueue.scala 154:109:@1693.4]
  assign _T_3542 = _T_3541 & noConflicts_7; // @[StoreQueue.scala 154:109:@1694.4]
  assign _T_3543 = _T_3542 & noConflicts_8; // @[StoreQueue.scala 154:109:@1695.4]
  assign _T_3544 = _T_3543 & noConflicts_9; // @[StoreQueue.scala 154:109:@1696.4]
  assign _T_3545 = _T_3544 & noConflicts_10; // @[StoreQueue.scala 154:109:@1697.4]
  assign _T_3546 = _T_3545 & noConflicts_11; // @[StoreQueue.scala 154:109:@1698.4]
  assign _T_3547 = _T_3546 & noConflicts_12; // @[StoreQueue.scala 154:109:@1699.4]
  assign _T_3548 = _T_3547 & noConflicts_13; // @[StoreQueue.scala 154:109:@1700.4]
  assign _T_3549 = _T_3548 & noConflicts_14; // @[StoreQueue.scala 154:109:@1701.4]
  assign _T_3550 = _T_3549 & noConflicts_15; // @[StoreQueue.scala 154:109:@1702.4]
  assign storeRequest = _T_3533 & _T_3550; // @[StoreQueue.scala 154:88:@1703.4]
  assign _T_3553 = head == 4'h0; // @[StoreQueue.scala 164:23:@1708.6]
  assign _T_3554 = _T_3553 & storeRequest; // @[StoreQueue.scala 164:43:@1709.6]
  assign _T_3555 = _T_3554 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1710.6]
  assign _GEN_960 = _T_3555 ? 1'h1 : storeCompleted_0; // @[StoreQueue.scala 164:86:@1711.6]
  assign _GEN_961 = initBits_0 ? 1'h0 : _GEN_960; // @[StoreQueue.scala 162:37:@1704.4]
  assign _T_3559 = head == 4'h1; // @[StoreQueue.scala 164:23:@1718.6]
  assign _T_3560 = _T_3559 & storeRequest; // @[StoreQueue.scala 164:43:@1719.6]
  assign _T_3561 = _T_3560 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1720.6]
  assign _GEN_962 = _T_3561 ? 1'h1 : storeCompleted_1; // @[StoreQueue.scala 164:86:@1721.6]
  assign _GEN_963 = initBits_1 ? 1'h0 : _GEN_962; // @[StoreQueue.scala 162:37:@1714.4]
  assign _T_3565 = head == 4'h2; // @[StoreQueue.scala 164:23:@1728.6]
  assign _T_3566 = _T_3565 & storeRequest; // @[StoreQueue.scala 164:43:@1729.6]
  assign _T_3567 = _T_3566 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1730.6]
  assign _GEN_964 = _T_3567 ? 1'h1 : storeCompleted_2; // @[StoreQueue.scala 164:86:@1731.6]
  assign _GEN_965 = initBits_2 ? 1'h0 : _GEN_964; // @[StoreQueue.scala 162:37:@1724.4]
  assign _T_3571 = head == 4'h3; // @[StoreQueue.scala 164:23:@1738.6]
  assign _T_3572 = _T_3571 & storeRequest; // @[StoreQueue.scala 164:43:@1739.6]
  assign _T_3573 = _T_3572 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1740.6]
  assign _GEN_966 = _T_3573 ? 1'h1 : storeCompleted_3; // @[StoreQueue.scala 164:86:@1741.6]
  assign _GEN_967 = initBits_3 ? 1'h0 : _GEN_966; // @[StoreQueue.scala 162:37:@1734.4]
  assign _T_3577 = head == 4'h4; // @[StoreQueue.scala 164:23:@1748.6]
  assign _T_3578 = _T_3577 & storeRequest; // @[StoreQueue.scala 164:43:@1749.6]
  assign _T_3579 = _T_3578 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1750.6]
  assign _GEN_968 = _T_3579 ? 1'h1 : storeCompleted_4; // @[StoreQueue.scala 164:86:@1751.6]
  assign _GEN_969 = initBits_4 ? 1'h0 : _GEN_968; // @[StoreQueue.scala 162:37:@1744.4]
  assign _T_3583 = head == 4'h5; // @[StoreQueue.scala 164:23:@1758.6]
  assign _T_3584 = _T_3583 & storeRequest; // @[StoreQueue.scala 164:43:@1759.6]
  assign _T_3585 = _T_3584 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1760.6]
  assign _GEN_970 = _T_3585 ? 1'h1 : storeCompleted_5; // @[StoreQueue.scala 164:86:@1761.6]
  assign _GEN_971 = initBits_5 ? 1'h0 : _GEN_970; // @[StoreQueue.scala 162:37:@1754.4]
  assign _T_3589 = head == 4'h6; // @[StoreQueue.scala 164:23:@1768.6]
  assign _T_3590 = _T_3589 & storeRequest; // @[StoreQueue.scala 164:43:@1769.6]
  assign _T_3591 = _T_3590 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1770.6]
  assign _GEN_972 = _T_3591 ? 1'h1 : storeCompleted_6; // @[StoreQueue.scala 164:86:@1771.6]
  assign _GEN_973 = initBits_6 ? 1'h0 : _GEN_972; // @[StoreQueue.scala 162:37:@1764.4]
  assign _T_3595 = head == 4'h7; // @[StoreQueue.scala 164:23:@1778.6]
  assign _T_3596 = _T_3595 & storeRequest; // @[StoreQueue.scala 164:43:@1779.6]
  assign _T_3597 = _T_3596 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1780.6]
  assign _GEN_974 = _T_3597 ? 1'h1 : storeCompleted_7; // @[StoreQueue.scala 164:86:@1781.6]
  assign _GEN_975 = initBits_7 ? 1'h0 : _GEN_974; // @[StoreQueue.scala 162:37:@1774.4]
  assign _T_3601 = head == 4'h8; // @[StoreQueue.scala 164:23:@1788.6]
  assign _T_3602 = _T_3601 & storeRequest; // @[StoreQueue.scala 164:43:@1789.6]
  assign _T_3603 = _T_3602 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1790.6]
  assign _GEN_976 = _T_3603 ? 1'h1 : storeCompleted_8; // @[StoreQueue.scala 164:86:@1791.6]
  assign _GEN_977 = initBits_8 ? 1'h0 : _GEN_976; // @[StoreQueue.scala 162:37:@1784.4]
  assign _T_3607 = head == 4'h9; // @[StoreQueue.scala 164:23:@1798.6]
  assign _T_3608 = _T_3607 & storeRequest; // @[StoreQueue.scala 164:43:@1799.6]
  assign _T_3609 = _T_3608 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1800.6]
  assign _GEN_978 = _T_3609 ? 1'h1 : storeCompleted_9; // @[StoreQueue.scala 164:86:@1801.6]
  assign _GEN_979 = initBits_9 ? 1'h0 : _GEN_978; // @[StoreQueue.scala 162:37:@1794.4]
  assign _T_3613 = head == 4'ha; // @[StoreQueue.scala 164:23:@1808.6]
  assign _T_3614 = _T_3613 & storeRequest; // @[StoreQueue.scala 164:43:@1809.6]
  assign _T_3615 = _T_3614 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1810.6]
  assign _GEN_980 = _T_3615 ? 1'h1 : storeCompleted_10; // @[StoreQueue.scala 164:86:@1811.6]
  assign _GEN_981 = initBits_10 ? 1'h0 : _GEN_980; // @[StoreQueue.scala 162:37:@1804.4]
  assign _T_3619 = head == 4'hb; // @[StoreQueue.scala 164:23:@1818.6]
  assign _T_3620 = _T_3619 & storeRequest; // @[StoreQueue.scala 164:43:@1819.6]
  assign _T_3621 = _T_3620 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1820.6]
  assign _GEN_982 = _T_3621 ? 1'h1 : storeCompleted_11; // @[StoreQueue.scala 164:86:@1821.6]
  assign _GEN_983 = initBits_11 ? 1'h0 : _GEN_982; // @[StoreQueue.scala 162:37:@1814.4]
  assign _T_3625 = head == 4'hc; // @[StoreQueue.scala 164:23:@1828.6]
  assign _T_3626 = _T_3625 & storeRequest; // @[StoreQueue.scala 164:43:@1829.6]
  assign _T_3627 = _T_3626 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1830.6]
  assign _GEN_984 = _T_3627 ? 1'h1 : storeCompleted_12; // @[StoreQueue.scala 164:86:@1831.6]
  assign _GEN_985 = initBits_12 ? 1'h0 : _GEN_984; // @[StoreQueue.scala 162:37:@1824.4]
  assign _T_3631 = head == 4'hd; // @[StoreQueue.scala 164:23:@1838.6]
  assign _T_3632 = _T_3631 & storeRequest; // @[StoreQueue.scala 164:43:@1839.6]
  assign _T_3633 = _T_3632 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1840.6]
  assign _GEN_986 = _T_3633 ? 1'h1 : storeCompleted_13; // @[StoreQueue.scala 164:86:@1841.6]
  assign _GEN_987 = initBits_13 ? 1'h0 : _GEN_986; // @[StoreQueue.scala 162:37:@1834.4]
  assign _T_3637 = head == 4'he; // @[StoreQueue.scala 164:23:@1848.6]
  assign _T_3638 = _T_3637 & storeRequest; // @[StoreQueue.scala 164:43:@1849.6]
  assign _T_3639 = _T_3638 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1850.6]
  assign _GEN_988 = _T_3639 ? 1'h1 : storeCompleted_14; // @[StoreQueue.scala 164:86:@1851.6]
  assign _GEN_989 = initBits_14 ? 1'h0 : _GEN_988; // @[StoreQueue.scala 162:37:@1844.4]
  assign _T_3643 = head == 4'hf; // @[StoreQueue.scala 164:23:@1858.6]
  assign _T_3644 = _T_3643 & storeRequest; // @[StoreQueue.scala 164:43:@1859.6]
  assign _T_3645 = _T_3644 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1860.6]
  assign _GEN_990 = _T_3645 ? 1'h1 : storeCompleted_15; // @[StoreQueue.scala 164:86:@1861.6]
  assign _GEN_991 = initBits_15 ? 1'h0 : _GEN_990; // @[StoreQueue.scala 162:37:@1854.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[StoreQueue.scala 180:72:@1865.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[StoreQueue.scala 180:72:@1867.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[StoreQueue.scala 180:72:@1869.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[StoreQueue.scala 180:72:@1871.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[StoreQueue.scala 180:72:@1873.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[StoreQueue.scala 180:72:@1875.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[StoreQueue.scala 180:72:@1877.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[StoreQueue.scala 180:72:@1879.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[StoreQueue.scala 180:72:@1881.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[StoreQueue.scala 180:72:@1883.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[StoreQueue.scala 180:72:@1885.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[StoreQueue.scala 180:72:@1887.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[StoreQueue.scala 180:72:@1889.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[StoreQueue.scala 180:72:@1891.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[StoreQueue.scala 180:72:@1893.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[StoreQueue.scala 180:72:@1895.4]
  assign _T_4378 = addrKnown_0 == 1'h0; // @[StoreQueue.scala 192:91:@1931.4]
  assign _T_4379 = entriesPorts_0_0 & _T_4378; // @[StoreQueue.scala 192:88:@1932.4]
  assign _T_4381 = addrKnown_1 == 1'h0; // @[StoreQueue.scala 192:91:@1933.4]
  assign _T_4382 = entriesPorts_0_1 & _T_4381; // @[StoreQueue.scala 192:88:@1934.4]
  assign _T_4384 = addrKnown_2 == 1'h0; // @[StoreQueue.scala 192:91:@1935.4]
  assign _T_4385 = entriesPorts_0_2 & _T_4384; // @[StoreQueue.scala 192:88:@1936.4]
  assign _T_4387 = addrKnown_3 == 1'h0; // @[StoreQueue.scala 192:91:@1937.4]
  assign _T_4388 = entriesPorts_0_3 & _T_4387; // @[StoreQueue.scala 192:88:@1938.4]
  assign _T_4390 = addrKnown_4 == 1'h0; // @[StoreQueue.scala 192:91:@1939.4]
  assign _T_4391 = entriesPorts_0_4 & _T_4390; // @[StoreQueue.scala 192:88:@1940.4]
  assign _T_4393 = addrKnown_5 == 1'h0; // @[StoreQueue.scala 192:91:@1941.4]
  assign _T_4394 = entriesPorts_0_5 & _T_4393; // @[StoreQueue.scala 192:88:@1942.4]
  assign _T_4396 = addrKnown_6 == 1'h0; // @[StoreQueue.scala 192:91:@1943.4]
  assign _T_4397 = entriesPorts_0_6 & _T_4396; // @[StoreQueue.scala 192:88:@1944.4]
  assign _T_4399 = addrKnown_7 == 1'h0; // @[StoreQueue.scala 192:91:@1945.4]
  assign _T_4400 = entriesPorts_0_7 & _T_4399; // @[StoreQueue.scala 192:88:@1946.4]
  assign _T_4402 = addrKnown_8 == 1'h0; // @[StoreQueue.scala 192:91:@1947.4]
  assign _T_4403 = entriesPorts_0_8 & _T_4402; // @[StoreQueue.scala 192:88:@1948.4]
  assign _T_4405 = addrKnown_9 == 1'h0; // @[StoreQueue.scala 192:91:@1949.4]
  assign _T_4406 = entriesPorts_0_9 & _T_4405; // @[StoreQueue.scala 192:88:@1950.4]
  assign _T_4408 = addrKnown_10 == 1'h0; // @[StoreQueue.scala 192:91:@1951.4]
  assign _T_4409 = entriesPorts_0_10 & _T_4408; // @[StoreQueue.scala 192:88:@1952.4]
  assign _T_4411 = addrKnown_11 == 1'h0; // @[StoreQueue.scala 192:91:@1953.4]
  assign _T_4412 = entriesPorts_0_11 & _T_4411; // @[StoreQueue.scala 192:88:@1954.4]
  assign _T_4414 = addrKnown_12 == 1'h0; // @[StoreQueue.scala 192:91:@1955.4]
  assign _T_4415 = entriesPorts_0_12 & _T_4414; // @[StoreQueue.scala 192:88:@1956.4]
  assign _T_4417 = addrKnown_13 == 1'h0; // @[StoreQueue.scala 192:91:@1957.4]
  assign _T_4418 = entriesPorts_0_13 & _T_4417; // @[StoreQueue.scala 192:88:@1958.4]
  assign _T_4420 = addrKnown_14 == 1'h0; // @[StoreQueue.scala 192:91:@1959.4]
  assign _T_4421 = entriesPorts_0_14 & _T_4420; // @[StoreQueue.scala 192:88:@1960.4]
  assign _T_4423 = addrKnown_15 == 1'h0; // @[StoreQueue.scala 192:91:@1961.4]
  assign _T_4424 = entriesPorts_0_15 & _T_4423; // @[StoreQueue.scala 192:88:@1962.4]
  assign _T_4448 = dataKnown_0 == 1'h0; // @[StoreQueue.scala 193:91:@1980.4]
  assign _T_4449 = entriesPorts_0_0 & _T_4448; // @[StoreQueue.scala 193:88:@1981.4]
  assign _T_4451 = dataKnown_1 == 1'h0; // @[StoreQueue.scala 193:91:@1982.4]
  assign _T_4452 = entriesPorts_0_1 & _T_4451; // @[StoreQueue.scala 193:88:@1983.4]
  assign _T_4454 = dataKnown_2 == 1'h0; // @[StoreQueue.scala 193:91:@1984.4]
  assign _T_4455 = entriesPorts_0_2 & _T_4454; // @[StoreQueue.scala 193:88:@1985.4]
  assign _T_4457 = dataKnown_3 == 1'h0; // @[StoreQueue.scala 193:91:@1986.4]
  assign _T_4458 = entriesPorts_0_3 & _T_4457; // @[StoreQueue.scala 193:88:@1987.4]
  assign _T_4460 = dataKnown_4 == 1'h0; // @[StoreQueue.scala 193:91:@1988.4]
  assign _T_4461 = entriesPorts_0_4 & _T_4460; // @[StoreQueue.scala 193:88:@1989.4]
  assign _T_4463 = dataKnown_5 == 1'h0; // @[StoreQueue.scala 193:91:@1990.4]
  assign _T_4464 = entriesPorts_0_5 & _T_4463; // @[StoreQueue.scala 193:88:@1991.4]
  assign _T_4466 = dataKnown_6 == 1'h0; // @[StoreQueue.scala 193:91:@1992.4]
  assign _T_4467 = entriesPorts_0_6 & _T_4466; // @[StoreQueue.scala 193:88:@1993.4]
  assign _T_4469 = dataKnown_7 == 1'h0; // @[StoreQueue.scala 193:91:@1994.4]
  assign _T_4470 = entriesPorts_0_7 & _T_4469; // @[StoreQueue.scala 193:88:@1995.4]
  assign _T_4472 = dataKnown_8 == 1'h0; // @[StoreQueue.scala 193:91:@1996.4]
  assign _T_4473 = entriesPorts_0_8 & _T_4472; // @[StoreQueue.scala 193:88:@1997.4]
  assign _T_4475 = dataKnown_9 == 1'h0; // @[StoreQueue.scala 193:91:@1998.4]
  assign _T_4476 = entriesPorts_0_9 & _T_4475; // @[StoreQueue.scala 193:88:@1999.4]
  assign _T_4478 = dataKnown_10 == 1'h0; // @[StoreQueue.scala 193:91:@2000.4]
  assign _T_4479 = entriesPorts_0_10 & _T_4478; // @[StoreQueue.scala 193:88:@2001.4]
  assign _T_4481 = dataKnown_11 == 1'h0; // @[StoreQueue.scala 193:91:@2002.4]
  assign _T_4482 = entriesPorts_0_11 & _T_4481; // @[StoreQueue.scala 193:88:@2003.4]
  assign _T_4484 = dataKnown_12 == 1'h0; // @[StoreQueue.scala 193:91:@2004.4]
  assign _T_4485 = entriesPorts_0_12 & _T_4484; // @[StoreQueue.scala 193:88:@2005.4]
  assign _T_4487 = dataKnown_13 == 1'h0; // @[StoreQueue.scala 193:91:@2006.4]
  assign _T_4488 = entriesPorts_0_13 & _T_4487; // @[StoreQueue.scala 193:88:@2007.4]
  assign _T_4490 = dataKnown_14 == 1'h0; // @[StoreQueue.scala 193:91:@2008.4]
  assign _T_4491 = entriesPorts_0_14 & _T_4490; // @[StoreQueue.scala 193:88:@2009.4]
  assign _T_4493 = dataKnown_15 == 1'h0; // @[StoreQueue.scala 193:91:@2010.4]
  assign _T_4494 = entriesPorts_0_15 & _T_4493; // @[StoreQueue.scala 193:88:@2011.4]
  assign _T_4519 = 16'h1 << head; // @[OneHot.scala 52:12:@2030.4]
  assign _T_4521 = _T_4519[0]; // @[util.scala 33:60:@2032.4]
  assign _T_4522 = _T_4519[1]; // @[util.scala 33:60:@2033.4]
  assign _T_4523 = _T_4519[2]; // @[util.scala 33:60:@2034.4]
  assign _T_4524 = _T_4519[3]; // @[util.scala 33:60:@2035.4]
  assign _T_4525 = _T_4519[4]; // @[util.scala 33:60:@2036.4]
  assign _T_4526 = _T_4519[5]; // @[util.scala 33:60:@2037.4]
  assign _T_4527 = _T_4519[6]; // @[util.scala 33:60:@2038.4]
  assign _T_4528 = _T_4519[7]; // @[util.scala 33:60:@2039.4]
  assign _T_4529 = _T_4519[8]; // @[util.scala 33:60:@2040.4]
  assign _T_4530 = _T_4519[9]; // @[util.scala 33:60:@2041.4]
  assign _T_4531 = _T_4519[10]; // @[util.scala 33:60:@2042.4]
  assign _T_4532 = _T_4519[11]; // @[util.scala 33:60:@2043.4]
  assign _T_4533 = _T_4519[12]; // @[util.scala 33:60:@2044.4]
  assign _T_4534 = _T_4519[13]; // @[util.scala 33:60:@2045.4]
  assign _T_4535 = _T_4519[14]; // @[util.scala 33:60:@2046.4]
  assign _T_4536 = _T_4519[15]; // @[util.scala 33:60:@2047.4]
  assign _T_4577 = _T_4424 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2065.4]
  assign _T_4578 = _T_4421 ? 16'h4000 : _T_4577; // @[Mux.scala 31:69:@2066.4]
  assign _T_4579 = _T_4418 ? 16'h2000 : _T_4578; // @[Mux.scala 31:69:@2067.4]
  assign _T_4580 = _T_4415 ? 16'h1000 : _T_4579; // @[Mux.scala 31:69:@2068.4]
  assign _T_4581 = _T_4412 ? 16'h800 : _T_4580; // @[Mux.scala 31:69:@2069.4]
  assign _T_4582 = _T_4409 ? 16'h400 : _T_4581; // @[Mux.scala 31:69:@2070.4]
  assign _T_4583 = _T_4406 ? 16'h200 : _T_4582; // @[Mux.scala 31:69:@2071.4]
  assign _T_4584 = _T_4403 ? 16'h100 : _T_4583; // @[Mux.scala 31:69:@2072.4]
  assign _T_4585 = _T_4400 ? 16'h80 : _T_4584; // @[Mux.scala 31:69:@2073.4]
  assign _T_4586 = _T_4397 ? 16'h40 : _T_4585; // @[Mux.scala 31:69:@2074.4]
  assign _T_4587 = _T_4394 ? 16'h20 : _T_4586; // @[Mux.scala 31:69:@2075.4]
  assign _T_4588 = _T_4391 ? 16'h10 : _T_4587; // @[Mux.scala 31:69:@2076.4]
  assign _T_4589 = _T_4388 ? 16'h8 : _T_4588; // @[Mux.scala 31:69:@2077.4]
  assign _T_4590 = _T_4385 ? 16'h4 : _T_4589; // @[Mux.scala 31:69:@2078.4]
  assign _T_4591 = _T_4382 ? 16'h2 : _T_4590; // @[Mux.scala 31:69:@2079.4]
  assign _T_4592 = _T_4379 ? 16'h1 : _T_4591; // @[Mux.scala 31:69:@2080.4]
  assign _T_4593 = _T_4592[0]; // @[OneHot.scala 66:30:@2081.4]
  assign _T_4594 = _T_4592[1]; // @[OneHot.scala 66:30:@2082.4]
  assign _T_4595 = _T_4592[2]; // @[OneHot.scala 66:30:@2083.4]
  assign _T_4596 = _T_4592[3]; // @[OneHot.scala 66:30:@2084.4]
  assign _T_4597 = _T_4592[4]; // @[OneHot.scala 66:30:@2085.4]
  assign _T_4598 = _T_4592[5]; // @[OneHot.scala 66:30:@2086.4]
  assign _T_4599 = _T_4592[6]; // @[OneHot.scala 66:30:@2087.4]
  assign _T_4600 = _T_4592[7]; // @[OneHot.scala 66:30:@2088.4]
  assign _T_4601 = _T_4592[8]; // @[OneHot.scala 66:30:@2089.4]
  assign _T_4602 = _T_4592[9]; // @[OneHot.scala 66:30:@2090.4]
  assign _T_4603 = _T_4592[10]; // @[OneHot.scala 66:30:@2091.4]
  assign _T_4604 = _T_4592[11]; // @[OneHot.scala 66:30:@2092.4]
  assign _T_4605 = _T_4592[12]; // @[OneHot.scala 66:30:@2093.4]
  assign _T_4606 = _T_4592[13]; // @[OneHot.scala 66:30:@2094.4]
  assign _T_4607 = _T_4592[14]; // @[OneHot.scala 66:30:@2095.4]
  assign _T_4608 = _T_4592[15]; // @[OneHot.scala 66:30:@2096.4]
  assign _T_4649 = _T_4379 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2114.4]
  assign _T_4650 = _T_4424 ? 16'h4000 : _T_4649; // @[Mux.scala 31:69:@2115.4]
  assign _T_4651 = _T_4421 ? 16'h2000 : _T_4650; // @[Mux.scala 31:69:@2116.4]
  assign _T_4652 = _T_4418 ? 16'h1000 : _T_4651; // @[Mux.scala 31:69:@2117.4]
  assign _T_4653 = _T_4415 ? 16'h800 : _T_4652; // @[Mux.scala 31:69:@2118.4]
  assign _T_4654 = _T_4412 ? 16'h400 : _T_4653; // @[Mux.scala 31:69:@2119.4]
  assign _T_4655 = _T_4409 ? 16'h200 : _T_4654; // @[Mux.scala 31:69:@2120.4]
  assign _T_4656 = _T_4406 ? 16'h100 : _T_4655; // @[Mux.scala 31:69:@2121.4]
  assign _T_4657 = _T_4403 ? 16'h80 : _T_4656; // @[Mux.scala 31:69:@2122.4]
  assign _T_4658 = _T_4400 ? 16'h40 : _T_4657; // @[Mux.scala 31:69:@2123.4]
  assign _T_4659 = _T_4397 ? 16'h20 : _T_4658; // @[Mux.scala 31:69:@2124.4]
  assign _T_4660 = _T_4394 ? 16'h10 : _T_4659; // @[Mux.scala 31:69:@2125.4]
  assign _T_4661 = _T_4391 ? 16'h8 : _T_4660; // @[Mux.scala 31:69:@2126.4]
  assign _T_4662 = _T_4388 ? 16'h4 : _T_4661; // @[Mux.scala 31:69:@2127.4]
  assign _T_4663 = _T_4385 ? 16'h2 : _T_4662; // @[Mux.scala 31:69:@2128.4]
  assign _T_4664 = _T_4382 ? 16'h1 : _T_4663; // @[Mux.scala 31:69:@2129.4]
  assign _T_4665 = _T_4664[0]; // @[OneHot.scala 66:30:@2130.4]
  assign _T_4666 = _T_4664[1]; // @[OneHot.scala 66:30:@2131.4]
  assign _T_4667 = _T_4664[2]; // @[OneHot.scala 66:30:@2132.4]
  assign _T_4668 = _T_4664[3]; // @[OneHot.scala 66:30:@2133.4]
  assign _T_4669 = _T_4664[4]; // @[OneHot.scala 66:30:@2134.4]
  assign _T_4670 = _T_4664[5]; // @[OneHot.scala 66:30:@2135.4]
  assign _T_4671 = _T_4664[6]; // @[OneHot.scala 66:30:@2136.4]
  assign _T_4672 = _T_4664[7]; // @[OneHot.scala 66:30:@2137.4]
  assign _T_4673 = _T_4664[8]; // @[OneHot.scala 66:30:@2138.4]
  assign _T_4674 = _T_4664[9]; // @[OneHot.scala 66:30:@2139.4]
  assign _T_4675 = _T_4664[10]; // @[OneHot.scala 66:30:@2140.4]
  assign _T_4676 = _T_4664[11]; // @[OneHot.scala 66:30:@2141.4]
  assign _T_4677 = _T_4664[12]; // @[OneHot.scala 66:30:@2142.4]
  assign _T_4678 = _T_4664[13]; // @[OneHot.scala 66:30:@2143.4]
  assign _T_4679 = _T_4664[14]; // @[OneHot.scala 66:30:@2144.4]
  assign _T_4680 = _T_4664[15]; // @[OneHot.scala 66:30:@2145.4]
  assign _T_4721 = _T_4382 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2163.4]
  assign _T_4722 = _T_4379 ? 16'h4000 : _T_4721; // @[Mux.scala 31:69:@2164.4]
  assign _T_4723 = _T_4424 ? 16'h2000 : _T_4722; // @[Mux.scala 31:69:@2165.4]
  assign _T_4724 = _T_4421 ? 16'h1000 : _T_4723; // @[Mux.scala 31:69:@2166.4]
  assign _T_4725 = _T_4418 ? 16'h800 : _T_4724; // @[Mux.scala 31:69:@2167.4]
  assign _T_4726 = _T_4415 ? 16'h400 : _T_4725; // @[Mux.scala 31:69:@2168.4]
  assign _T_4727 = _T_4412 ? 16'h200 : _T_4726; // @[Mux.scala 31:69:@2169.4]
  assign _T_4728 = _T_4409 ? 16'h100 : _T_4727; // @[Mux.scala 31:69:@2170.4]
  assign _T_4729 = _T_4406 ? 16'h80 : _T_4728; // @[Mux.scala 31:69:@2171.4]
  assign _T_4730 = _T_4403 ? 16'h40 : _T_4729; // @[Mux.scala 31:69:@2172.4]
  assign _T_4731 = _T_4400 ? 16'h20 : _T_4730; // @[Mux.scala 31:69:@2173.4]
  assign _T_4732 = _T_4397 ? 16'h10 : _T_4731; // @[Mux.scala 31:69:@2174.4]
  assign _T_4733 = _T_4394 ? 16'h8 : _T_4732; // @[Mux.scala 31:69:@2175.4]
  assign _T_4734 = _T_4391 ? 16'h4 : _T_4733; // @[Mux.scala 31:69:@2176.4]
  assign _T_4735 = _T_4388 ? 16'h2 : _T_4734; // @[Mux.scala 31:69:@2177.4]
  assign _T_4736 = _T_4385 ? 16'h1 : _T_4735; // @[Mux.scala 31:69:@2178.4]
  assign _T_4737 = _T_4736[0]; // @[OneHot.scala 66:30:@2179.4]
  assign _T_4738 = _T_4736[1]; // @[OneHot.scala 66:30:@2180.4]
  assign _T_4739 = _T_4736[2]; // @[OneHot.scala 66:30:@2181.4]
  assign _T_4740 = _T_4736[3]; // @[OneHot.scala 66:30:@2182.4]
  assign _T_4741 = _T_4736[4]; // @[OneHot.scala 66:30:@2183.4]
  assign _T_4742 = _T_4736[5]; // @[OneHot.scala 66:30:@2184.4]
  assign _T_4743 = _T_4736[6]; // @[OneHot.scala 66:30:@2185.4]
  assign _T_4744 = _T_4736[7]; // @[OneHot.scala 66:30:@2186.4]
  assign _T_4745 = _T_4736[8]; // @[OneHot.scala 66:30:@2187.4]
  assign _T_4746 = _T_4736[9]; // @[OneHot.scala 66:30:@2188.4]
  assign _T_4747 = _T_4736[10]; // @[OneHot.scala 66:30:@2189.4]
  assign _T_4748 = _T_4736[11]; // @[OneHot.scala 66:30:@2190.4]
  assign _T_4749 = _T_4736[12]; // @[OneHot.scala 66:30:@2191.4]
  assign _T_4750 = _T_4736[13]; // @[OneHot.scala 66:30:@2192.4]
  assign _T_4751 = _T_4736[14]; // @[OneHot.scala 66:30:@2193.4]
  assign _T_4752 = _T_4736[15]; // @[OneHot.scala 66:30:@2194.4]
  assign _T_4793 = _T_4385 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2212.4]
  assign _T_4794 = _T_4382 ? 16'h4000 : _T_4793; // @[Mux.scala 31:69:@2213.4]
  assign _T_4795 = _T_4379 ? 16'h2000 : _T_4794; // @[Mux.scala 31:69:@2214.4]
  assign _T_4796 = _T_4424 ? 16'h1000 : _T_4795; // @[Mux.scala 31:69:@2215.4]
  assign _T_4797 = _T_4421 ? 16'h800 : _T_4796; // @[Mux.scala 31:69:@2216.4]
  assign _T_4798 = _T_4418 ? 16'h400 : _T_4797; // @[Mux.scala 31:69:@2217.4]
  assign _T_4799 = _T_4415 ? 16'h200 : _T_4798; // @[Mux.scala 31:69:@2218.4]
  assign _T_4800 = _T_4412 ? 16'h100 : _T_4799; // @[Mux.scala 31:69:@2219.4]
  assign _T_4801 = _T_4409 ? 16'h80 : _T_4800; // @[Mux.scala 31:69:@2220.4]
  assign _T_4802 = _T_4406 ? 16'h40 : _T_4801; // @[Mux.scala 31:69:@2221.4]
  assign _T_4803 = _T_4403 ? 16'h20 : _T_4802; // @[Mux.scala 31:69:@2222.4]
  assign _T_4804 = _T_4400 ? 16'h10 : _T_4803; // @[Mux.scala 31:69:@2223.4]
  assign _T_4805 = _T_4397 ? 16'h8 : _T_4804; // @[Mux.scala 31:69:@2224.4]
  assign _T_4806 = _T_4394 ? 16'h4 : _T_4805; // @[Mux.scala 31:69:@2225.4]
  assign _T_4807 = _T_4391 ? 16'h2 : _T_4806; // @[Mux.scala 31:69:@2226.4]
  assign _T_4808 = _T_4388 ? 16'h1 : _T_4807; // @[Mux.scala 31:69:@2227.4]
  assign _T_4809 = _T_4808[0]; // @[OneHot.scala 66:30:@2228.4]
  assign _T_4810 = _T_4808[1]; // @[OneHot.scala 66:30:@2229.4]
  assign _T_4811 = _T_4808[2]; // @[OneHot.scala 66:30:@2230.4]
  assign _T_4812 = _T_4808[3]; // @[OneHot.scala 66:30:@2231.4]
  assign _T_4813 = _T_4808[4]; // @[OneHot.scala 66:30:@2232.4]
  assign _T_4814 = _T_4808[5]; // @[OneHot.scala 66:30:@2233.4]
  assign _T_4815 = _T_4808[6]; // @[OneHot.scala 66:30:@2234.4]
  assign _T_4816 = _T_4808[7]; // @[OneHot.scala 66:30:@2235.4]
  assign _T_4817 = _T_4808[8]; // @[OneHot.scala 66:30:@2236.4]
  assign _T_4818 = _T_4808[9]; // @[OneHot.scala 66:30:@2237.4]
  assign _T_4819 = _T_4808[10]; // @[OneHot.scala 66:30:@2238.4]
  assign _T_4820 = _T_4808[11]; // @[OneHot.scala 66:30:@2239.4]
  assign _T_4821 = _T_4808[12]; // @[OneHot.scala 66:30:@2240.4]
  assign _T_4822 = _T_4808[13]; // @[OneHot.scala 66:30:@2241.4]
  assign _T_4823 = _T_4808[14]; // @[OneHot.scala 66:30:@2242.4]
  assign _T_4824 = _T_4808[15]; // @[OneHot.scala 66:30:@2243.4]
  assign _T_4865 = _T_4388 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2261.4]
  assign _T_4866 = _T_4385 ? 16'h4000 : _T_4865; // @[Mux.scala 31:69:@2262.4]
  assign _T_4867 = _T_4382 ? 16'h2000 : _T_4866; // @[Mux.scala 31:69:@2263.4]
  assign _T_4868 = _T_4379 ? 16'h1000 : _T_4867; // @[Mux.scala 31:69:@2264.4]
  assign _T_4869 = _T_4424 ? 16'h800 : _T_4868; // @[Mux.scala 31:69:@2265.4]
  assign _T_4870 = _T_4421 ? 16'h400 : _T_4869; // @[Mux.scala 31:69:@2266.4]
  assign _T_4871 = _T_4418 ? 16'h200 : _T_4870; // @[Mux.scala 31:69:@2267.4]
  assign _T_4872 = _T_4415 ? 16'h100 : _T_4871; // @[Mux.scala 31:69:@2268.4]
  assign _T_4873 = _T_4412 ? 16'h80 : _T_4872; // @[Mux.scala 31:69:@2269.4]
  assign _T_4874 = _T_4409 ? 16'h40 : _T_4873; // @[Mux.scala 31:69:@2270.4]
  assign _T_4875 = _T_4406 ? 16'h20 : _T_4874; // @[Mux.scala 31:69:@2271.4]
  assign _T_4876 = _T_4403 ? 16'h10 : _T_4875; // @[Mux.scala 31:69:@2272.4]
  assign _T_4877 = _T_4400 ? 16'h8 : _T_4876; // @[Mux.scala 31:69:@2273.4]
  assign _T_4878 = _T_4397 ? 16'h4 : _T_4877; // @[Mux.scala 31:69:@2274.4]
  assign _T_4879 = _T_4394 ? 16'h2 : _T_4878; // @[Mux.scala 31:69:@2275.4]
  assign _T_4880 = _T_4391 ? 16'h1 : _T_4879; // @[Mux.scala 31:69:@2276.4]
  assign _T_4881 = _T_4880[0]; // @[OneHot.scala 66:30:@2277.4]
  assign _T_4882 = _T_4880[1]; // @[OneHot.scala 66:30:@2278.4]
  assign _T_4883 = _T_4880[2]; // @[OneHot.scala 66:30:@2279.4]
  assign _T_4884 = _T_4880[3]; // @[OneHot.scala 66:30:@2280.4]
  assign _T_4885 = _T_4880[4]; // @[OneHot.scala 66:30:@2281.4]
  assign _T_4886 = _T_4880[5]; // @[OneHot.scala 66:30:@2282.4]
  assign _T_4887 = _T_4880[6]; // @[OneHot.scala 66:30:@2283.4]
  assign _T_4888 = _T_4880[7]; // @[OneHot.scala 66:30:@2284.4]
  assign _T_4889 = _T_4880[8]; // @[OneHot.scala 66:30:@2285.4]
  assign _T_4890 = _T_4880[9]; // @[OneHot.scala 66:30:@2286.4]
  assign _T_4891 = _T_4880[10]; // @[OneHot.scala 66:30:@2287.4]
  assign _T_4892 = _T_4880[11]; // @[OneHot.scala 66:30:@2288.4]
  assign _T_4893 = _T_4880[12]; // @[OneHot.scala 66:30:@2289.4]
  assign _T_4894 = _T_4880[13]; // @[OneHot.scala 66:30:@2290.4]
  assign _T_4895 = _T_4880[14]; // @[OneHot.scala 66:30:@2291.4]
  assign _T_4896 = _T_4880[15]; // @[OneHot.scala 66:30:@2292.4]
  assign _T_4937 = _T_4391 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2310.4]
  assign _T_4938 = _T_4388 ? 16'h4000 : _T_4937; // @[Mux.scala 31:69:@2311.4]
  assign _T_4939 = _T_4385 ? 16'h2000 : _T_4938; // @[Mux.scala 31:69:@2312.4]
  assign _T_4940 = _T_4382 ? 16'h1000 : _T_4939; // @[Mux.scala 31:69:@2313.4]
  assign _T_4941 = _T_4379 ? 16'h800 : _T_4940; // @[Mux.scala 31:69:@2314.4]
  assign _T_4942 = _T_4424 ? 16'h400 : _T_4941; // @[Mux.scala 31:69:@2315.4]
  assign _T_4943 = _T_4421 ? 16'h200 : _T_4942; // @[Mux.scala 31:69:@2316.4]
  assign _T_4944 = _T_4418 ? 16'h100 : _T_4943; // @[Mux.scala 31:69:@2317.4]
  assign _T_4945 = _T_4415 ? 16'h80 : _T_4944; // @[Mux.scala 31:69:@2318.4]
  assign _T_4946 = _T_4412 ? 16'h40 : _T_4945; // @[Mux.scala 31:69:@2319.4]
  assign _T_4947 = _T_4409 ? 16'h20 : _T_4946; // @[Mux.scala 31:69:@2320.4]
  assign _T_4948 = _T_4406 ? 16'h10 : _T_4947; // @[Mux.scala 31:69:@2321.4]
  assign _T_4949 = _T_4403 ? 16'h8 : _T_4948; // @[Mux.scala 31:69:@2322.4]
  assign _T_4950 = _T_4400 ? 16'h4 : _T_4949; // @[Mux.scala 31:69:@2323.4]
  assign _T_4951 = _T_4397 ? 16'h2 : _T_4950; // @[Mux.scala 31:69:@2324.4]
  assign _T_4952 = _T_4394 ? 16'h1 : _T_4951; // @[Mux.scala 31:69:@2325.4]
  assign _T_4953 = _T_4952[0]; // @[OneHot.scala 66:30:@2326.4]
  assign _T_4954 = _T_4952[1]; // @[OneHot.scala 66:30:@2327.4]
  assign _T_4955 = _T_4952[2]; // @[OneHot.scala 66:30:@2328.4]
  assign _T_4956 = _T_4952[3]; // @[OneHot.scala 66:30:@2329.4]
  assign _T_4957 = _T_4952[4]; // @[OneHot.scala 66:30:@2330.4]
  assign _T_4958 = _T_4952[5]; // @[OneHot.scala 66:30:@2331.4]
  assign _T_4959 = _T_4952[6]; // @[OneHot.scala 66:30:@2332.4]
  assign _T_4960 = _T_4952[7]; // @[OneHot.scala 66:30:@2333.4]
  assign _T_4961 = _T_4952[8]; // @[OneHot.scala 66:30:@2334.4]
  assign _T_4962 = _T_4952[9]; // @[OneHot.scala 66:30:@2335.4]
  assign _T_4963 = _T_4952[10]; // @[OneHot.scala 66:30:@2336.4]
  assign _T_4964 = _T_4952[11]; // @[OneHot.scala 66:30:@2337.4]
  assign _T_4965 = _T_4952[12]; // @[OneHot.scala 66:30:@2338.4]
  assign _T_4966 = _T_4952[13]; // @[OneHot.scala 66:30:@2339.4]
  assign _T_4967 = _T_4952[14]; // @[OneHot.scala 66:30:@2340.4]
  assign _T_4968 = _T_4952[15]; // @[OneHot.scala 66:30:@2341.4]
  assign _T_5009 = _T_4394 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2359.4]
  assign _T_5010 = _T_4391 ? 16'h4000 : _T_5009; // @[Mux.scala 31:69:@2360.4]
  assign _T_5011 = _T_4388 ? 16'h2000 : _T_5010; // @[Mux.scala 31:69:@2361.4]
  assign _T_5012 = _T_4385 ? 16'h1000 : _T_5011; // @[Mux.scala 31:69:@2362.4]
  assign _T_5013 = _T_4382 ? 16'h800 : _T_5012; // @[Mux.scala 31:69:@2363.4]
  assign _T_5014 = _T_4379 ? 16'h400 : _T_5013; // @[Mux.scala 31:69:@2364.4]
  assign _T_5015 = _T_4424 ? 16'h200 : _T_5014; // @[Mux.scala 31:69:@2365.4]
  assign _T_5016 = _T_4421 ? 16'h100 : _T_5015; // @[Mux.scala 31:69:@2366.4]
  assign _T_5017 = _T_4418 ? 16'h80 : _T_5016; // @[Mux.scala 31:69:@2367.4]
  assign _T_5018 = _T_4415 ? 16'h40 : _T_5017; // @[Mux.scala 31:69:@2368.4]
  assign _T_5019 = _T_4412 ? 16'h20 : _T_5018; // @[Mux.scala 31:69:@2369.4]
  assign _T_5020 = _T_4409 ? 16'h10 : _T_5019; // @[Mux.scala 31:69:@2370.4]
  assign _T_5021 = _T_4406 ? 16'h8 : _T_5020; // @[Mux.scala 31:69:@2371.4]
  assign _T_5022 = _T_4403 ? 16'h4 : _T_5021; // @[Mux.scala 31:69:@2372.4]
  assign _T_5023 = _T_4400 ? 16'h2 : _T_5022; // @[Mux.scala 31:69:@2373.4]
  assign _T_5024 = _T_4397 ? 16'h1 : _T_5023; // @[Mux.scala 31:69:@2374.4]
  assign _T_5025 = _T_5024[0]; // @[OneHot.scala 66:30:@2375.4]
  assign _T_5026 = _T_5024[1]; // @[OneHot.scala 66:30:@2376.4]
  assign _T_5027 = _T_5024[2]; // @[OneHot.scala 66:30:@2377.4]
  assign _T_5028 = _T_5024[3]; // @[OneHot.scala 66:30:@2378.4]
  assign _T_5029 = _T_5024[4]; // @[OneHot.scala 66:30:@2379.4]
  assign _T_5030 = _T_5024[5]; // @[OneHot.scala 66:30:@2380.4]
  assign _T_5031 = _T_5024[6]; // @[OneHot.scala 66:30:@2381.4]
  assign _T_5032 = _T_5024[7]; // @[OneHot.scala 66:30:@2382.4]
  assign _T_5033 = _T_5024[8]; // @[OneHot.scala 66:30:@2383.4]
  assign _T_5034 = _T_5024[9]; // @[OneHot.scala 66:30:@2384.4]
  assign _T_5035 = _T_5024[10]; // @[OneHot.scala 66:30:@2385.4]
  assign _T_5036 = _T_5024[11]; // @[OneHot.scala 66:30:@2386.4]
  assign _T_5037 = _T_5024[12]; // @[OneHot.scala 66:30:@2387.4]
  assign _T_5038 = _T_5024[13]; // @[OneHot.scala 66:30:@2388.4]
  assign _T_5039 = _T_5024[14]; // @[OneHot.scala 66:30:@2389.4]
  assign _T_5040 = _T_5024[15]; // @[OneHot.scala 66:30:@2390.4]
  assign _T_5081 = _T_4397 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2408.4]
  assign _T_5082 = _T_4394 ? 16'h4000 : _T_5081; // @[Mux.scala 31:69:@2409.4]
  assign _T_5083 = _T_4391 ? 16'h2000 : _T_5082; // @[Mux.scala 31:69:@2410.4]
  assign _T_5084 = _T_4388 ? 16'h1000 : _T_5083; // @[Mux.scala 31:69:@2411.4]
  assign _T_5085 = _T_4385 ? 16'h800 : _T_5084; // @[Mux.scala 31:69:@2412.4]
  assign _T_5086 = _T_4382 ? 16'h400 : _T_5085; // @[Mux.scala 31:69:@2413.4]
  assign _T_5087 = _T_4379 ? 16'h200 : _T_5086; // @[Mux.scala 31:69:@2414.4]
  assign _T_5088 = _T_4424 ? 16'h100 : _T_5087; // @[Mux.scala 31:69:@2415.4]
  assign _T_5089 = _T_4421 ? 16'h80 : _T_5088; // @[Mux.scala 31:69:@2416.4]
  assign _T_5090 = _T_4418 ? 16'h40 : _T_5089; // @[Mux.scala 31:69:@2417.4]
  assign _T_5091 = _T_4415 ? 16'h20 : _T_5090; // @[Mux.scala 31:69:@2418.4]
  assign _T_5092 = _T_4412 ? 16'h10 : _T_5091; // @[Mux.scala 31:69:@2419.4]
  assign _T_5093 = _T_4409 ? 16'h8 : _T_5092; // @[Mux.scala 31:69:@2420.4]
  assign _T_5094 = _T_4406 ? 16'h4 : _T_5093; // @[Mux.scala 31:69:@2421.4]
  assign _T_5095 = _T_4403 ? 16'h2 : _T_5094; // @[Mux.scala 31:69:@2422.4]
  assign _T_5096 = _T_4400 ? 16'h1 : _T_5095; // @[Mux.scala 31:69:@2423.4]
  assign _T_5097 = _T_5096[0]; // @[OneHot.scala 66:30:@2424.4]
  assign _T_5098 = _T_5096[1]; // @[OneHot.scala 66:30:@2425.4]
  assign _T_5099 = _T_5096[2]; // @[OneHot.scala 66:30:@2426.4]
  assign _T_5100 = _T_5096[3]; // @[OneHot.scala 66:30:@2427.4]
  assign _T_5101 = _T_5096[4]; // @[OneHot.scala 66:30:@2428.4]
  assign _T_5102 = _T_5096[5]; // @[OneHot.scala 66:30:@2429.4]
  assign _T_5103 = _T_5096[6]; // @[OneHot.scala 66:30:@2430.4]
  assign _T_5104 = _T_5096[7]; // @[OneHot.scala 66:30:@2431.4]
  assign _T_5105 = _T_5096[8]; // @[OneHot.scala 66:30:@2432.4]
  assign _T_5106 = _T_5096[9]; // @[OneHot.scala 66:30:@2433.4]
  assign _T_5107 = _T_5096[10]; // @[OneHot.scala 66:30:@2434.4]
  assign _T_5108 = _T_5096[11]; // @[OneHot.scala 66:30:@2435.4]
  assign _T_5109 = _T_5096[12]; // @[OneHot.scala 66:30:@2436.4]
  assign _T_5110 = _T_5096[13]; // @[OneHot.scala 66:30:@2437.4]
  assign _T_5111 = _T_5096[14]; // @[OneHot.scala 66:30:@2438.4]
  assign _T_5112 = _T_5096[15]; // @[OneHot.scala 66:30:@2439.4]
  assign _T_5153 = _T_4400 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2457.4]
  assign _T_5154 = _T_4397 ? 16'h4000 : _T_5153; // @[Mux.scala 31:69:@2458.4]
  assign _T_5155 = _T_4394 ? 16'h2000 : _T_5154; // @[Mux.scala 31:69:@2459.4]
  assign _T_5156 = _T_4391 ? 16'h1000 : _T_5155; // @[Mux.scala 31:69:@2460.4]
  assign _T_5157 = _T_4388 ? 16'h800 : _T_5156; // @[Mux.scala 31:69:@2461.4]
  assign _T_5158 = _T_4385 ? 16'h400 : _T_5157; // @[Mux.scala 31:69:@2462.4]
  assign _T_5159 = _T_4382 ? 16'h200 : _T_5158; // @[Mux.scala 31:69:@2463.4]
  assign _T_5160 = _T_4379 ? 16'h100 : _T_5159; // @[Mux.scala 31:69:@2464.4]
  assign _T_5161 = _T_4424 ? 16'h80 : _T_5160; // @[Mux.scala 31:69:@2465.4]
  assign _T_5162 = _T_4421 ? 16'h40 : _T_5161; // @[Mux.scala 31:69:@2466.4]
  assign _T_5163 = _T_4418 ? 16'h20 : _T_5162; // @[Mux.scala 31:69:@2467.4]
  assign _T_5164 = _T_4415 ? 16'h10 : _T_5163; // @[Mux.scala 31:69:@2468.4]
  assign _T_5165 = _T_4412 ? 16'h8 : _T_5164; // @[Mux.scala 31:69:@2469.4]
  assign _T_5166 = _T_4409 ? 16'h4 : _T_5165; // @[Mux.scala 31:69:@2470.4]
  assign _T_5167 = _T_4406 ? 16'h2 : _T_5166; // @[Mux.scala 31:69:@2471.4]
  assign _T_5168 = _T_4403 ? 16'h1 : _T_5167; // @[Mux.scala 31:69:@2472.4]
  assign _T_5169 = _T_5168[0]; // @[OneHot.scala 66:30:@2473.4]
  assign _T_5170 = _T_5168[1]; // @[OneHot.scala 66:30:@2474.4]
  assign _T_5171 = _T_5168[2]; // @[OneHot.scala 66:30:@2475.4]
  assign _T_5172 = _T_5168[3]; // @[OneHot.scala 66:30:@2476.4]
  assign _T_5173 = _T_5168[4]; // @[OneHot.scala 66:30:@2477.4]
  assign _T_5174 = _T_5168[5]; // @[OneHot.scala 66:30:@2478.4]
  assign _T_5175 = _T_5168[6]; // @[OneHot.scala 66:30:@2479.4]
  assign _T_5176 = _T_5168[7]; // @[OneHot.scala 66:30:@2480.4]
  assign _T_5177 = _T_5168[8]; // @[OneHot.scala 66:30:@2481.4]
  assign _T_5178 = _T_5168[9]; // @[OneHot.scala 66:30:@2482.4]
  assign _T_5179 = _T_5168[10]; // @[OneHot.scala 66:30:@2483.4]
  assign _T_5180 = _T_5168[11]; // @[OneHot.scala 66:30:@2484.4]
  assign _T_5181 = _T_5168[12]; // @[OneHot.scala 66:30:@2485.4]
  assign _T_5182 = _T_5168[13]; // @[OneHot.scala 66:30:@2486.4]
  assign _T_5183 = _T_5168[14]; // @[OneHot.scala 66:30:@2487.4]
  assign _T_5184 = _T_5168[15]; // @[OneHot.scala 66:30:@2488.4]
  assign _T_5225 = _T_4403 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2506.4]
  assign _T_5226 = _T_4400 ? 16'h4000 : _T_5225; // @[Mux.scala 31:69:@2507.4]
  assign _T_5227 = _T_4397 ? 16'h2000 : _T_5226; // @[Mux.scala 31:69:@2508.4]
  assign _T_5228 = _T_4394 ? 16'h1000 : _T_5227; // @[Mux.scala 31:69:@2509.4]
  assign _T_5229 = _T_4391 ? 16'h800 : _T_5228; // @[Mux.scala 31:69:@2510.4]
  assign _T_5230 = _T_4388 ? 16'h400 : _T_5229; // @[Mux.scala 31:69:@2511.4]
  assign _T_5231 = _T_4385 ? 16'h200 : _T_5230; // @[Mux.scala 31:69:@2512.4]
  assign _T_5232 = _T_4382 ? 16'h100 : _T_5231; // @[Mux.scala 31:69:@2513.4]
  assign _T_5233 = _T_4379 ? 16'h80 : _T_5232; // @[Mux.scala 31:69:@2514.4]
  assign _T_5234 = _T_4424 ? 16'h40 : _T_5233; // @[Mux.scala 31:69:@2515.4]
  assign _T_5235 = _T_4421 ? 16'h20 : _T_5234; // @[Mux.scala 31:69:@2516.4]
  assign _T_5236 = _T_4418 ? 16'h10 : _T_5235; // @[Mux.scala 31:69:@2517.4]
  assign _T_5237 = _T_4415 ? 16'h8 : _T_5236; // @[Mux.scala 31:69:@2518.4]
  assign _T_5238 = _T_4412 ? 16'h4 : _T_5237; // @[Mux.scala 31:69:@2519.4]
  assign _T_5239 = _T_4409 ? 16'h2 : _T_5238; // @[Mux.scala 31:69:@2520.4]
  assign _T_5240 = _T_4406 ? 16'h1 : _T_5239; // @[Mux.scala 31:69:@2521.4]
  assign _T_5241 = _T_5240[0]; // @[OneHot.scala 66:30:@2522.4]
  assign _T_5242 = _T_5240[1]; // @[OneHot.scala 66:30:@2523.4]
  assign _T_5243 = _T_5240[2]; // @[OneHot.scala 66:30:@2524.4]
  assign _T_5244 = _T_5240[3]; // @[OneHot.scala 66:30:@2525.4]
  assign _T_5245 = _T_5240[4]; // @[OneHot.scala 66:30:@2526.4]
  assign _T_5246 = _T_5240[5]; // @[OneHot.scala 66:30:@2527.4]
  assign _T_5247 = _T_5240[6]; // @[OneHot.scala 66:30:@2528.4]
  assign _T_5248 = _T_5240[7]; // @[OneHot.scala 66:30:@2529.4]
  assign _T_5249 = _T_5240[8]; // @[OneHot.scala 66:30:@2530.4]
  assign _T_5250 = _T_5240[9]; // @[OneHot.scala 66:30:@2531.4]
  assign _T_5251 = _T_5240[10]; // @[OneHot.scala 66:30:@2532.4]
  assign _T_5252 = _T_5240[11]; // @[OneHot.scala 66:30:@2533.4]
  assign _T_5253 = _T_5240[12]; // @[OneHot.scala 66:30:@2534.4]
  assign _T_5254 = _T_5240[13]; // @[OneHot.scala 66:30:@2535.4]
  assign _T_5255 = _T_5240[14]; // @[OneHot.scala 66:30:@2536.4]
  assign _T_5256 = _T_5240[15]; // @[OneHot.scala 66:30:@2537.4]
  assign _T_5297 = _T_4406 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2555.4]
  assign _T_5298 = _T_4403 ? 16'h4000 : _T_5297; // @[Mux.scala 31:69:@2556.4]
  assign _T_5299 = _T_4400 ? 16'h2000 : _T_5298; // @[Mux.scala 31:69:@2557.4]
  assign _T_5300 = _T_4397 ? 16'h1000 : _T_5299; // @[Mux.scala 31:69:@2558.4]
  assign _T_5301 = _T_4394 ? 16'h800 : _T_5300; // @[Mux.scala 31:69:@2559.4]
  assign _T_5302 = _T_4391 ? 16'h400 : _T_5301; // @[Mux.scala 31:69:@2560.4]
  assign _T_5303 = _T_4388 ? 16'h200 : _T_5302; // @[Mux.scala 31:69:@2561.4]
  assign _T_5304 = _T_4385 ? 16'h100 : _T_5303; // @[Mux.scala 31:69:@2562.4]
  assign _T_5305 = _T_4382 ? 16'h80 : _T_5304; // @[Mux.scala 31:69:@2563.4]
  assign _T_5306 = _T_4379 ? 16'h40 : _T_5305; // @[Mux.scala 31:69:@2564.4]
  assign _T_5307 = _T_4424 ? 16'h20 : _T_5306; // @[Mux.scala 31:69:@2565.4]
  assign _T_5308 = _T_4421 ? 16'h10 : _T_5307; // @[Mux.scala 31:69:@2566.4]
  assign _T_5309 = _T_4418 ? 16'h8 : _T_5308; // @[Mux.scala 31:69:@2567.4]
  assign _T_5310 = _T_4415 ? 16'h4 : _T_5309; // @[Mux.scala 31:69:@2568.4]
  assign _T_5311 = _T_4412 ? 16'h2 : _T_5310; // @[Mux.scala 31:69:@2569.4]
  assign _T_5312 = _T_4409 ? 16'h1 : _T_5311; // @[Mux.scala 31:69:@2570.4]
  assign _T_5313 = _T_5312[0]; // @[OneHot.scala 66:30:@2571.4]
  assign _T_5314 = _T_5312[1]; // @[OneHot.scala 66:30:@2572.4]
  assign _T_5315 = _T_5312[2]; // @[OneHot.scala 66:30:@2573.4]
  assign _T_5316 = _T_5312[3]; // @[OneHot.scala 66:30:@2574.4]
  assign _T_5317 = _T_5312[4]; // @[OneHot.scala 66:30:@2575.4]
  assign _T_5318 = _T_5312[5]; // @[OneHot.scala 66:30:@2576.4]
  assign _T_5319 = _T_5312[6]; // @[OneHot.scala 66:30:@2577.4]
  assign _T_5320 = _T_5312[7]; // @[OneHot.scala 66:30:@2578.4]
  assign _T_5321 = _T_5312[8]; // @[OneHot.scala 66:30:@2579.4]
  assign _T_5322 = _T_5312[9]; // @[OneHot.scala 66:30:@2580.4]
  assign _T_5323 = _T_5312[10]; // @[OneHot.scala 66:30:@2581.4]
  assign _T_5324 = _T_5312[11]; // @[OneHot.scala 66:30:@2582.4]
  assign _T_5325 = _T_5312[12]; // @[OneHot.scala 66:30:@2583.4]
  assign _T_5326 = _T_5312[13]; // @[OneHot.scala 66:30:@2584.4]
  assign _T_5327 = _T_5312[14]; // @[OneHot.scala 66:30:@2585.4]
  assign _T_5328 = _T_5312[15]; // @[OneHot.scala 66:30:@2586.4]
  assign _T_5369 = _T_4409 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2604.4]
  assign _T_5370 = _T_4406 ? 16'h4000 : _T_5369; // @[Mux.scala 31:69:@2605.4]
  assign _T_5371 = _T_4403 ? 16'h2000 : _T_5370; // @[Mux.scala 31:69:@2606.4]
  assign _T_5372 = _T_4400 ? 16'h1000 : _T_5371; // @[Mux.scala 31:69:@2607.4]
  assign _T_5373 = _T_4397 ? 16'h800 : _T_5372; // @[Mux.scala 31:69:@2608.4]
  assign _T_5374 = _T_4394 ? 16'h400 : _T_5373; // @[Mux.scala 31:69:@2609.4]
  assign _T_5375 = _T_4391 ? 16'h200 : _T_5374; // @[Mux.scala 31:69:@2610.4]
  assign _T_5376 = _T_4388 ? 16'h100 : _T_5375; // @[Mux.scala 31:69:@2611.4]
  assign _T_5377 = _T_4385 ? 16'h80 : _T_5376; // @[Mux.scala 31:69:@2612.4]
  assign _T_5378 = _T_4382 ? 16'h40 : _T_5377; // @[Mux.scala 31:69:@2613.4]
  assign _T_5379 = _T_4379 ? 16'h20 : _T_5378; // @[Mux.scala 31:69:@2614.4]
  assign _T_5380 = _T_4424 ? 16'h10 : _T_5379; // @[Mux.scala 31:69:@2615.4]
  assign _T_5381 = _T_4421 ? 16'h8 : _T_5380; // @[Mux.scala 31:69:@2616.4]
  assign _T_5382 = _T_4418 ? 16'h4 : _T_5381; // @[Mux.scala 31:69:@2617.4]
  assign _T_5383 = _T_4415 ? 16'h2 : _T_5382; // @[Mux.scala 31:69:@2618.4]
  assign _T_5384 = _T_4412 ? 16'h1 : _T_5383; // @[Mux.scala 31:69:@2619.4]
  assign _T_5385 = _T_5384[0]; // @[OneHot.scala 66:30:@2620.4]
  assign _T_5386 = _T_5384[1]; // @[OneHot.scala 66:30:@2621.4]
  assign _T_5387 = _T_5384[2]; // @[OneHot.scala 66:30:@2622.4]
  assign _T_5388 = _T_5384[3]; // @[OneHot.scala 66:30:@2623.4]
  assign _T_5389 = _T_5384[4]; // @[OneHot.scala 66:30:@2624.4]
  assign _T_5390 = _T_5384[5]; // @[OneHot.scala 66:30:@2625.4]
  assign _T_5391 = _T_5384[6]; // @[OneHot.scala 66:30:@2626.4]
  assign _T_5392 = _T_5384[7]; // @[OneHot.scala 66:30:@2627.4]
  assign _T_5393 = _T_5384[8]; // @[OneHot.scala 66:30:@2628.4]
  assign _T_5394 = _T_5384[9]; // @[OneHot.scala 66:30:@2629.4]
  assign _T_5395 = _T_5384[10]; // @[OneHot.scala 66:30:@2630.4]
  assign _T_5396 = _T_5384[11]; // @[OneHot.scala 66:30:@2631.4]
  assign _T_5397 = _T_5384[12]; // @[OneHot.scala 66:30:@2632.4]
  assign _T_5398 = _T_5384[13]; // @[OneHot.scala 66:30:@2633.4]
  assign _T_5399 = _T_5384[14]; // @[OneHot.scala 66:30:@2634.4]
  assign _T_5400 = _T_5384[15]; // @[OneHot.scala 66:30:@2635.4]
  assign _T_5441 = _T_4412 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2653.4]
  assign _T_5442 = _T_4409 ? 16'h4000 : _T_5441; // @[Mux.scala 31:69:@2654.4]
  assign _T_5443 = _T_4406 ? 16'h2000 : _T_5442; // @[Mux.scala 31:69:@2655.4]
  assign _T_5444 = _T_4403 ? 16'h1000 : _T_5443; // @[Mux.scala 31:69:@2656.4]
  assign _T_5445 = _T_4400 ? 16'h800 : _T_5444; // @[Mux.scala 31:69:@2657.4]
  assign _T_5446 = _T_4397 ? 16'h400 : _T_5445; // @[Mux.scala 31:69:@2658.4]
  assign _T_5447 = _T_4394 ? 16'h200 : _T_5446; // @[Mux.scala 31:69:@2659.4]
  assign _T_5448 = _T_4391 ? 16'h100 : _T_5447; // @[Mux.scala 31:69:@2660.4]
  assign _T_5449 = _T_4388 ? 16'h80 : _T_5448; // @[Mux.scala 31:69:@2661.4]
  assign _T_5450 = _T_4385 ? 16'h40 : _T_5449; // @[Mux.scala 31:69:@2662.4]
  assign _T_5451 = _T_4382 ? 16'h20 : _T_5450; // @[Mux.scala 31:69:@2663.4]
  assign _T_5452 = _T_4379 ? 16'h10 : _T_5451; // @[Mux.scala 31:69:@2664.4]
  assign _T_5453 = _T_4424 ? 16'h8 : _T_5452; // @[Mux.scala 31:69:@2665.4]
  assign _T_5454 = _T_4421 ? 16'h4 : _T_5453; // @[Mux.scala 31:69:@2666.4]
  assign _T_5455 = _T_4418 ? 16'h2 : _T_5454; // @[Mux.scala 31:69:@2667.4]
  assign _T_5456 = _T_4415 ? 16'h1 : _T_5455; // @[Mux.scala 31:69:@2668.4]
  assign _T_5457 = _T_5456[0]; // @[OneHot.scala 66:30:@2669.4]
  assign _T_5458 = _T_5456[1]; // @[OneHot.scala 66:30:@2670.4]
  assign _T_5459 = _T_5456[2]; // @[OneHot.scala 66:30:@2671.4]
  assign _T_5460 = _T_5456[3]; // @[OneHot.scala 66:30:@2672.4]
  assign _T_5461 = _T_5456[4]; // @[OneHot.scala 66:30:@2673.4]
  assign _T_5462 = _T_5456[5]; // @[OneHot.scala 66:30:@2674.4]
  assign _T_5463 = _T_5456[6]; // @[OneHot.scala 66:30:@2675.4]
  assign _T_5464 = _T_5456[7]; // @[OneHot.scala 66:30:@2676.4]
  assign _T_5465 = _T_5456[8]; // @[OneHot.scala 66:30:@2677.4]
  assign _T_5466 = _T_5456[9]; // @[OneHot.scala 66:30:@2678.4]
  assign _T_5467 = _T_5456[10]; // @[OneHot.scala 66:30:@2679.4]
  assign _T_5468 = _T_5456[11]; // @[OneHot.scala 66:30:@2680.4]
  assign _T_5469 = _T_5456[12]; // @[OneHot.scala 66:30:@2681.4]
  assign _T_5470 = _T_5456[13]; // @[OneHot.scala 66:30:@2682.4]
  assign _T_5471 = _T_5456[14]; // @[OneHot.scala 66:30:@2683.4]
  assign _T_5472 = _T_5456[15]; // @[OneHot.scala 66:30:@2684.4]
  assign _T_5513 = _T_4415 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2702.4]
  assign _T_5514 = _T_4412 ? 16'h4000 : _T_5513; // @[Mux.scala 31:69:@2703.4]
  assign _T_5515 = _T_4409 ? 16'h2000 : _T_5514; // @[Mux.scala 31:69:@2704.4]
  assign _T_5516 = _T_4406 ? 16'h1000 : _T_5515; // @[Mux.scala 31:69:@2705.4]
  assign _T_5517 = _T_4403 ? 16'h800 : _T_5516; // @[Mux.scala 31:69:@2706.4]
  assign _T_5518 = _T_4400 ? 16'h400 : _T_5517; // @[Mux.scala 31:69:@2707.4]
  assign _T_5519 = _T_4397 ? 16'h200 : _T_5518; // @[Mux.scala 31:69:@2708.4]
  assign _T_5520 = _T_4394 ? 16'h100 : _T_5519; // @[Mux.scala 31:69:@2709.4]
  assign _T_5521 = _T_4391 ? 16'h80 : _T_5520; // @[Mux.scala 31:69:@2710.4]
  assign _T_5522 = _T_4388 ? 16'h40 : _T_5521; // @[Mux.scala 31:69:@2711.4]
  assign _T_5523 = _T_4385 ? 16'h20 : _T_5522; // @[Mux.scala 31:69:@2712.4]
  assign _T_5524 = _T_4382 ? 16'h10 : _T_5523; // @[Mux.scala 31:69:@2713.4]
  assign _T_5525 = _T_4379 ? 16'h8 : _T_5524; // @[Mux.scala 31:69:@2714.4]
  assign _T_5526 = _T_4424 ? 16'h4 : _T_5525; // @[Mux.scala 31:69:@2715.4]
  assign _T_5527 = _T_4421 ? 16'h2 : _T_5526; // @[Mux.scala 31:69:@2716.4]
  assign _T_5528 = _T_4418 ? 16'h1 : _T_5527; // @[Mux.scala 31:69:@2717.4]
  assign _T_5529 = _T_5528[0]; // @[OneHot.scala 66:30:@2718.4]
  assign _T_5530 = _T_5528[1]; // @[OneHot.scala 66:30:@2719.4]
  assign _T_5531 = _T_5528[2]; // @[OneHot.scala 66:30:@2720.4]
  assign _T_5532 = _T_5528[3]; // @[OneHot.scala 66:30:@2721.4]
  assign _T_5533 = _T_5528[4]; // @[OneHot.scala 66:30:@2722.4]
  assign _T_5534 = _T_5528[5]; // @[OneHot.scala 66:30:@2723.4]
  assign _T_5535 = _T_5528[6]; // @[OneHot.scala 66:30:@2724.4]
  assign _T_5536 = _T_5528[7]; // @[OneHot.scala 66:30:@2725.4]
  assign _T_5537 = _T_5528[8]; // @[OneHot.scala 66:30:@2726.4]
  assign _T_5538 = _T_5528[9]; // @[OneHot.scala 66:30:@2727.4]
  assign _T_5539 = _T_5528[10]; // @[OneHot.scala 66:30:@2728.4]
  assign _T_5540 = _T_5528[11]; // @[OneHot.scala 66:30:@2729.4]
  assign _T_5541 = _T_5528[12]; // @[OneHot.scala 66:30:@2730.4]
  assign _T_5542 = _T_5528[13]; // @[OneHot.scala 66:30:@2731.4]
  assign _T_5543 = _T_5528[14]; // @[OneHot.scala 66:30:@2732.4]
  assign _T_5544 = _T_5528[15]; // @[OneHot.scala 66:30:@2733.4]
  assign _T_5585 = _T_4418 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2751.4]
  assign _T_5586 = _T_4415 ? 16'h4000 : _T_5585; // @[Mux.scala 31:69:@2752.4]
  assign _T_5587 = _T_4412 ? 16'h2000 : _T_5586; // @[Mux.scala 31:69:@2753.4]
  assign _T_5588 = _T_4409 ? 16'h1000 : _T_5587; // @[Mux.scala 31:69:@2754.4]
  assign _T_5589 = _T_4406 ? 16'h800 : _T_5588; // @[Mux.scala 31:69:@2755.4]
  assign _T_5590 = _T_4403 ? 16'h400 : _T_5589; // @[Mux.scala 31:69:@2756.4]
  assign _T_5591 = _T_4400 ? 16'h200 : _T_5590; // @[Mux.scala 31:69:@2757.4]
  assign _T_5592 = _T_4397 ? 16'h100 : _T_5591; // @[Mux.scala 31:69:@2758.4]
  assign _T_5593 = _T_4394 ? 16'h80 : _T_5592; // @[Mux.scala 31:69:@2759.4]
  assign _T_5594 = _T_4391 ? 16'h40 : _T_5593; // @[Mux.scala 31:69:@2760.4]
  assign _T_5595 = _T_4388 ? 16'h20 : _T_5594; // @[Mux.scala 31:69:@2761.4]
  assign _T_5596 = _T_4385 ? 16'h10 : _T_5595; // @[Mux.scala 31:69:@2762.4]
  assign _T_5597 = _T_4382 ? 16'h8 : _T_5596; // @[Mux.scala 31:69:@2763.4]
  assign _T_5598 = _T_4379 ? 16'h4 : _T_5597; // @[Mux.scala 31:69:@2764.4]
  assign _T_5599 = _T_4424 ? 16'h2 : _T_5598; // @[Mux.scala 31:69:@2765.4]
  assign _T_5600 = _T_4421 ? 16'h1 : _T_5599; // @[Mux.scala 31:69:@2766.4]
  assign _T_5601 = _T_5600[0]; // @[OneHot.scala 66:30:@2767.4]
  assign _T_5602 = _T_5600[1]; // @[OneHot.scala 66:30:@2768.4]
  assign _T_5603 = _T_5600[2]; // @[OneHot.scala 66:30:@2769.4]
  assign _T_5604 = _T_5600[3]; // @[OneHot.scala 66:30:@2770.4]
  assign _T_5605 = _T_5600[4]; // @[OneHot.scala 66:30:@2771.4]
  assign _T_5606 = _T_5600[5]; // @[OneHot.scala 66:30:@2772.4]
  assign _T_5607 = _T_5600[6]; // @[OneHot.scala 66:30:@2773.4]
  assign _T_5608 = _T_5600[7]; // @[OneHot.scala 66:30:@2774.4]
  assign _T_5609 = _T_5600[8]; // @[OneHot.scala 66:30:@2775.4]
  assign _T_5610 = _T_5600[9]; // @[OneHot.scala 66:30:@2776.4]
  assign _T_5611 = _T_5600[10]; // @[OneHot.scala 66:30:@2777.4]
  assign _T_5612 = _T_5600[11]; // @[OneHot.scala 66:30:@2778.4]
  assign _T_5613 = _T_5600[12]; // @[OneHot.scala 66:30:@2779.4]
  assign _T_5614 = _T_5600[13]; // @[OneHot.scala 66:30:@2780.4]
  assign _T_5615 = _T_5600[14]; // @[OneHot.scala 66:30:@2781.4]
  assign _T_5616 = _T_5600[15]; // @[OneHot.scala 66:30:@2782.4]
  assign _T_5657 = _T_4421 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2800.4]
  assign _T_5658 = _T_4418 ? 16'h4000 : _T_5657; // @[Mux.scala 31:69:@2801.4]
  assign _T_5659 = _T_4415 ? 16'h2000 : _T_5658; // @[Mux.scala 31:69:@2802.4]
  assign _T_5660 = _T_4412 ? 16'h1000 : _T_5659; // @[Mux.scala 31:69:@2803.4]
  assign _T_5661 = _T_4409 ? 16'h800 : _T_5660; // @[Mux.scala 31:69:@2804.4]
  assign _T_5662 = _T_4406 ? 16'h400 : _T_5661; // @[Mux.scala 31:69:@2805.4]
  assign _T_5663 = _T_4403 ? 16'h200 : _T_5662; // @[Mux.scala 31:69:@2806.4]
  assign _T_5664 = _T_4400 ? 16'h100 : _T_5663; // @[Mux.scala 31:69:@2807.4]
  assign _T_5665 = _T_4397 ? 16'h80 : _T_5664; // @[Mux.scala 31:69:@2808.4]
  assign _T_5666 = _T_4394 ? 16'h40 : _T_5665; // @[Mux.scala 31:69:@2809.4]
  assign _T_5667 = _T_4391 ? 16'h20 : _T_5666; // @[Mux.scala 31:69:@2810.4]
  assign _T_5668 = _T_4388 ? 16'h10 : _T_5667; // @[Mux.scala 31:69:@2811.4]
  assign _T_5669 = _T_4385 ? 16'h8 : _T_5668; // @[Mux.scala 31:69:@2812.4]
  assign _T_5670 = _T_4382 ? 16'h4 : _T_5669; // @[Mux.scala 31:69:@2813.4]
  assign _T_5671 = _T_4379 ? 16'h2 : _T_5670; // @[Mux.scala 31:69:@2814.4]
  assign _T_5672 = _T_4424 ? 16'h1 : _T_5671; // @[Mux.scala 31:69:@2815.4]
  assign _T_5673 = _T_5672[0]; // @[OneHot.scala 66:30:@2816.4]
  assign _T_5674 = _T_5672[1]; // @[OneHot.scala 66:30:@2817.4]
  assign _T_5675 = _T_5672[2]; // @[OneHot.scala 66:30:@2818.4]
  assign _T_5676 = _T_5672[3]; // @[OneHot.scala 66:30:@2819.4]
  assign _T_5677 = _T_5672[4]; // @[OneHot.scala 66:30:@2820.4]
  assign _T_5678 = _T_5672[5]; // @[OneHot.scala 66:30:@2821.4]
  assign _T_5679 = _T_5672[6]; // @[OneHot.scala 66:30:@2822.4]
  assign _T_5680 = _T_5672[7]; // @[OneHot.scala 66:30:@2823.4]
  assign _T_5681 = _T_5672[8]; // @[OneHot.scala 66:30:@2824.4]
  assign _T_5682 = _T_5672[9]; // @[OneHot.scala 66:30:@2825.4]
  assign _T_5683 = _T_5672[10]; // @[OneHot.scala 66:30:@2826.4]
  assign _T_5684 = _T_5672[11]; // @[OneHot.scala 66:30:@2827.4]
  assign _T_5685 = _T_5672[12]; // @[OneHot.scala 66:30:@2828.4]
  assign _T_5686 = _T_5672[13]; // @[OneHot.scala 66:30:@2829.4]
  assign _T_5687 = _T_5672[14]; // @[OneHot.scala 66:30:@2830.4]
  assign _T_5688 = _T_5672[15]; // @[OneHot.scala 66:30:@2831.4]
  assign _T_5753 = {_T_4600,_T_4599,_T_4598,_T_4597,_T_4596,_T_4595,_T_4594,_T_4593}; // @[Mux.scala 19:72:@2855.4]
  assign _T_5761 = {_T_4608,_T_4607,_T_4606,_T_4605,_T_4604,_T_4603,_T_4602,_T_4601,_T_5753}; // @[Mux.scala 19:72:@2863.4]
  assign _T_5763 = _T_4521 ? _T_5761 : 16'h0; // @[Mux.scala 19:72:@2864.4]
  assign _T_5770 = {_T_4671,_T_4670,_T_4669,_T_4668,_T_4667,_T_4666,_T_4665,_T_4680}; // @[Mux.scala 19:72:@2871.4]
  assign _T_5778 = {_T_4679,_T_4678,_T_4677,_T_4676,_T_4675,_T_4674,_T_4673,_T_4672,_T_5770}; // @[Mux.scala 19:72:@2879.4]
  assign _T_5780 = _T_4522 ? _T_5778 : 16'h0; // @[Mux.scala 19:72:@2880.4]
  assign _T_5787 = {_T_4742,_T_4741,_T_4740,_T_4739,_T_4738,_T_4737,_T_4752,_T_4751}; // @[Mux.scala 19:72:@2887.4]
  assign _T_5795 = {_T_4750,_T_4749,_T_4748,_T_4747,_T_4746,_T_4745,_T_4744,_T_4743,_T_5787}; // @[Mux.scala 19:72:@2895.4]
  assign _T_5797 = _T_4523 ? _T_5795 : 16'h0; // @[Mux.scala 19:72:@2896.4]
  assign _T_5804 = {_T_4813,_T_4812,_T_4811,_T_4810,_T_4809,_T_4824,_T_4823,_T_4822}; // @[Mux.scala 19:72:@2903.4]
  assign _T_5812 = {_T_4821,_T_4820,_T_4819,_T_4818,_T_4817,_T_4816,_T_4815,_T_4814,_T_5804}; // @[Mux.scala 19:72:@2911.4]
  assign _T_5814 = _T_4524 ? _T_5812 : 16'h0; // @[Mux.scala 19:72:@2912.4]
  assign _T_5821 = {_T_4884,_T_4883,_T_4882,_T_4881,_T_4896,_T_4895,_T_4894,_T_4893}; // @[Mux.scala 19:72:@2919.4]
  assign _T_5829 = {_T_4892,_T_4891,_T_4890,_T_4889,_T_4888,_T_4887,_T_4886,_T_4885,_T_5821}; // @[Mux.scala 19:72:@2927.4]
  assign _T_5831 = _T_4525 ? _T_5829 : 16'h0; // @[Mux.scala 19:72:@2928.4]
  assign _T_5838 = {_T_4955,_T_4954,_T_4953,_T_4968,_T_4967,_T_4966,_T_4965,_T_4964}; // @[Mux.scala 19:72:@2935.4]
  assign _T_5846 = {_T_4963,_T_4962,_T_4961,_T_4960,_T_4959,_T_4958,_T_4957,_T_4956,_T_5838}; // @[Mux.scala 19:72:@2943.4]
  assign _T_5848 = _T_4526 ? _T_5846 : 16'h0; // @[Mux.scala 19:72:@2944.4]
  assign _T_5855 = {_T_5026,_T_5025,_T_5040,_T_5039,_T_5038,_T_5037,_T_5036,_T_5035}; // @[Mux.scala 19:72:@2951.4]
  assign _T_5863 = {_T_5034,_T_5033,_T_5032,_T_5031,_T_5030,_T_5029,_T_5028,_T_5027,_T_5855}; // @[Mux.scala 19:72:@2959.4]
  assign _T_5865 = _T_4527 ? _T_5863 : 16'h0; // @[Mux.scala 19:72:@2960.4]
  assign _T_5872 = {_T_5097,_T_5112,_T_5111,_T_5110,_T_5109,_T_5108,_T_5107,_T_5106}; // @[Mux.scala 19:72:@2967.4]
  assign _T_5880 = {_T_5105,_T_5104,_T_5103,_T_5102,_T_5101,_T_5100,_T_5099,_T_5098,_T_5872}; // @[Mux.scala 19:72:@2975.4]
  assign _T_5882 = _T_4528 ? _T_5880 : 16'h0; // @[Mux.scala 19:72:@2976.4]
  assign _T_5889 = {_T_5184,_T_5183,_T_5182,_T_5181,_T_5180,_T_5179,_T_5178,_T_5177}; // @[Mux.scala 19:72:@2983.4]
  assign _T_5897 = {_T_5176,_T_5175,_T_5174,_T_5173,_T_5172,_T_5171,_T_5170,_T_5169,_T_5889}; // @[Mux.scala 19:72:@2991.4]
  assign _T_5899 = _T_4529 ? _T_5897 : 16'h0; // @[Mux.scala 19:72:@2992.4]
  assign _T_5906 = {_T_5255,_T_5254,_T_5253,_T_5252,_T_5251,_T_5250,_T_5249,_T_5248}; // @[Mux.scala 19:72:@2999.4]
  assign _T_5914 = {_T_5247,_T_5246,_T_5245,_T_5244,_T_5243,_T_5242,_T_5241,_T_5256,_T_5906}; // @[Mux.scala 19:72:@3007.4]
  assign _T_5916 = _T_4530 ? _T_5914 : 16'h0; // @[Mux.scala 19:72:@3008.4]
  assign _T_5923 = {_T_5326,_T_5325,_T_5324,_T_5323,_T_5322,_T_5321,_T_5320,_T_5319}; // @[Mux.scala 19:72:@3015.4]
  assign _T_5931 = {_T_5318,_T_5317,_T_5316,_T_5315,_T_5314,_T_5313,_T_5328,_T_5327,_T_5923}; // @[Mux.scala 19:72:@3023.4]
  assign _T_5933 = _T_4531 ? _T_5931 : 16'h0; // @[Mux.scala 19:72:@3024.4]
  assign _T_5940 = {_T_5397,_T_5396,_T_5395,_T_5394,_T_5393,_T_5392,_T_5391,_T_5390}; // @[Mux.scala 19:72:@3031.4]
  assign _T_5948 = {_T_5389,_T_5388,_T_5387,_T_5386,_T_5385,_T_5400,_T_5399,_T_5398,_T_5940}; // @[Mux.scala 19:72:@3039.4]
  assign _T_5950 = _T_4532 ? _T_5948 : 16'h0; // @[Mux.scala 19:72:@3040.4]
  assign _T_5957 = {_T_5468,_T_5467,_T_5466,_T_5465,_T_5464,_T_5463,_T_5462,_T_5461}; // @[Mux.scala 19:72:@3047.4]
  assign _T_5965 = {_T_5460,_T_5459,_T_5458,_T_5457,_T_5472,_T_5471,_T_5470,_T_5469,_T_5957}; // @[Mux.scala 19:72:@3055.4]
  assign _T_5967 = _T_4533 ? _T_5965 : 16'h0; // @[Mux.scala 19:72:@3056.4]
  assign _T_5974 = {_T_5539,_T_5538,_T_5537,_T_5536,_T_5535,_T_5534,_T_5533,_T_5532}; // @[Mux.scala 19:72:@3063.4]
  assign _T_5982 = {_T_5531,_T_5530,_T_5529,_T_5544,_T_5543,_T_5542,_T_5541,_T_5540,_T_5974}; // @[Mux.scala 19:72:@3071.4]
  assign _T_5984 = _T_4534 ? _T_5982 : 16'h0; // @[Mux.scala 19:72:@3072.4]
  assign _T_5991 = {_T_5610,_T_5609,_T_5608,_T_5607,_T_5606,_T_5605,_T_5604,_T_5603}; // @[Mux.scala 19:72:@3079.4]
  assign _T_5999 = {_T_5602,_T_5601,_T_5616,_T_5615,_T_5614,_T_5613,_T_5612,_T_5611,_T_5991}; // @[Mux.scala 19:72:@3087.4]
  assign _T_6001 = _T_4535 ? _T_5999 : 16'h0; // @[Mux.scala 19:72:@3088.4]
  assign _T_6008 = {_T_5681,_T_5680,_T_5679,_T_5678,_T_5677,_T_5676,_T_5675,_T_5674}; // @[Mux.scala 19:72:@3095.4]
  assign _T_6016 = {_T_5673,_T_5688,_T_5687,_T_5686,_T_5685,_T_5684,_T_5683,_T_5682,_T_6008}; // @[Mux.scala 19:72:@3103.4]
  assign _T_6018 = _T_4536 ? _T_6016 : 16'h0; // @[Mux.scala 19:72:@3104.4]
  assign _T_6019 = _T_5763 | _T_5780; // @[Mux.scala 19:72:@3105.4]
  assign _T_6020 = _T_6019 | _T_5797; // @[Mux.scala 19:72:@3106.4]
  assign _T_6021 = _T_6020 | _T_5814; // @[Mux.scala 19:72:@3107.4]
  assign _T_6022 = _T_6021 | _T_5831; // @[Mux.scala 19:72:@3108.4]
  assign _T_6023 = _T_6022 | _T_5848; // @[Mux.scala 19:72:@3109.4]
  assign _T_6024 = _T_6023 | _T_5865; // @[Mux.scala 19:72:@3110.4]
  assign _T_6025 = _T_6024 | _T_5882; // @[Mux.scala 19:72:@3111.4]
  assign _T_6026 = _T_6025 | _T_5899; // @[Mux.scala 19:72:@3112.4]
  assign _T_6027 = _T_6026 | _T_5916; // @[Mux.scala 19:72:@3113.4]
  assign _T_6028 = _T_6027 | _T_5933; // @[Mux.scala 19:72:@3114.4]
  assign _T_6029 = _T_6028 | _T_5950; // @[Mux.scala 19:72:@3115.4]
  assign _T_6030 = _T_6029 | _T_5967; // @[Mux.scala 19:72:@3116.4]
  assign _T_6031 = _T_6030 | _T_5984; // @[Mux.scala 19:72:@3117.4]
  assign _T_6032 = _T_6031 | _T_6001; // @[Mux.scala 19:72:@3118.4]
  assign _T_6033 = _T_6032 | _T_6018; // @[Mux.scala 19:72:@3119.4]
  assign inputAddrPriorityPorts_0_0 = _T_6033[0]; // @[Mux.scala 19:72:@3123.4]
  assign inputAddrPriorityPorts_0_1 = _T_6033[1]; // @[Mux.scala 19:72:@3125.4]
  assign inputAddrPriorityPorts_0_2 = _T_6033[2]; // @[Mux.scala 19:72:@3127.4]
  assign inputAddrPriorityPorts_0_3 = _T_6033[3]; // @[Mux.scala 19:72:@3129.4]
  assign inputAddrPriorityPorts_0_4 = _T_6033[4]; // @[Mux.scala 19:72:@3131.4]
  assign inputAddrPriorityPorts_0_5 = _T_6033[5]; // @[Mux.scala 19:72:@3133.4]
  assign inputAddrPriorityPorts_0_6 = _T_6033[6]; // @[Mux.scala 19:72:@3135.4]
  assign inputAddrPriorityPorts_0_7 = _T_6033[7]; // @[Mux.scala 19:72:@3137.4]
  assign inputAddrPriorityPorts_0_8 = _T_6033[8]; // @[Mux.scala 19:72:@3139.4]
  assign inputAddrPriorityPorts_0_9 = _T_6033[9]; // @[Mux.scala 19:72:@3141.4]
  assign inputAddrPriorityPorts_0_10 = _T_6033[10]; // @[Mux.scala 19:72:@3143.4]
  assign inputAddrPriorityPorts_0_11 = _T_6033[11]; // @[Mux.scala 19:72:@3145.4]
  assign inputAddrPriorityPorts_0_12 = _T_6033[12]; // @[Mux.scala 19:72:@3147.4]
  assign inputAddrPriorityPorts_0_13 = _T_6033[13]; // @[Mux.scala 19:72:@3149.4]
  assign inputAddrPriorityPorts_0_14 = _T_6033[14]; // @[Mux.scala 19:72:@3151.4]
  assign inputAddrPriorityPorts_0_15 = _T_6033[15]; // @[Mux.scala 19:72:@3153.4]
  assign _T_6235 = _T_4494 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3207.4]
  assign _T_6236 = _T_4491 ? 16'h4000 : _T_6235; // @[Mux.scala 31:69:@3208.4]
  assign _T_6237 = _T_4488 ? 16'h2000 : _T_6236; // @[Mux.scala 31:69:@3209.4]
  assign _T_6238 = _T_4485 ? 16'h1000 : _T_6237; // @[Mux.scala 31:69:@3210.4]
  assign _T_6239 = _T_4482 ? 16'h800 : _T_6238; // @[Mux.scala 31:69:@3211.4]
  assign _T_6240 = _T_4479 ? 16'h400 : _T_6239; // @[Mux.scala 31:69:@3212.4]
  assign _T_6241 = _T_4476 ? 16'h200 : _T_6240; // @[Mux.scala 31:69:@3213.4]
  assign _T_6242 = _T_4473 ? 16'h100 : _T_6241; // @[Mux.scala 31:69:@3214.4]
  assign _T_6243 = _T_4470 ? 16'h80 : _T_6242; // @[Mux.scala 31:69:@3215.4]
  assign _T_6244 = _T_4467 ? 16'h40 : _T_6243; // @[Mux.scala 31:69:@3216.4]
  assign _T_6245 = _T_4464 ? 16'h20 : _T_6244; // @[Mux.scala 31:69:@3217.4]
  assign _T_6246 = _T_4461 ? 16'h10 : _T_6245; // @[Mux.scala 31:69:@3218.4]
  assign _T_6247 = _T_4458 ? 16'h8 : _T_6246; // @[Mux.scala 31:69:@3219.4]
  assign _T_6248 = _T_4455 ? 16'h4 : _T_6247; // @[Mux.scala 31:69:@3220.4]
  assign _T_6249 = _T_4452 ? 16'h2 : _T_6248; // @[Mux.scala 31:69:@3221.4]
  assign _T_6250 = _T_4449 ? 16'h1 : _T_6249; // @[Mux.scala 31:69:@3222.4]
  assign _T_6251 = _T_6250[0]; // @[OneHot.scala 66:30:@3223.4]
  assign _T_6252 = _T_6250[1]; // @[OneHot.scala 66:30:@3224.4]
  assign _T_6253 = _T_6250[2]; // @[OneHot.scala 66:30:@3225.4]
  assign _T_6254 = _T_6250[3]; // @[OneHot.scala 66:30:@3226.4]
  assign _T_6255 = _T_6250[4]; // @[OneHot.scala 66:30:@3227.4]
  assign _T_6256 = _T_6250[5]; // @[OneHot.scala 66:30:@3228.4]
  assign _T_6257 = _T_6250[6]; // @[OneHot.scala 66:30:@3229.4]
  assign _T_6258 = _T_6250[7]; // @[OneHot.scala 66:30:@3230.4]
  assign _T_6259 = _T_6250[8]; // @[OneHot.scala 66:30:@3231.4]
  assign _T_6260 = _T_6250[9]; // @[OneHot.scala 66:30:@3232.4]
  assign _T_6261 = _T_6250[10]; // @[OneHot.scala 66:30:@3233.4]
  assign _T_6262 = _T_6250[11]; // @[OneHot.scala 66:30:@3234.4]
  assign _T_6263 = _T_6250[12]; // @[OneHot.scala 66:30:@3235.4]
  assign _T_6264 = _T_6250[13]; // @[OneHot.scala 66:30:@3236.4]
  assign _T_6265 = _T_6250[14]; // @[OneHot.scala 66:30:@3237.4]
  assign _T_6266 = _T_6250[15]; // @[OneHot.scala 66:30:@3238.4]
  assign _T_6307 = _T_4449 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3256.4]
  assign _T_6308 = _T_4494 ? 16'h4000 : _T_6307; // @[Mux.scala 31:69:@3257.4]
  assign _T_6309 = _T_4491 ? 16'h2000 : _T_6308; // @[Mux.scala 31:69:@3258.4]
  assign _T_6310 = _T_4488 ? 16'h1000 : _T_6309; // @[Mux.scala 31:69:@3259.4]
  assign _T_6311 = _T_4485 ? 16'h800 : _T_6310; // @[Mux.scala 31:69:@3260.4]
  assign _T_6312 = _T_4482 ? 16'h400 : _T_6311; // @[Mux.scala 31:69:@3261.4]
  assign _T_6313 = _T_4479 ? 16'h200 : _T_6312; // @[Mux.scala 31:69:@3262.4]
  assign _T_6314 = _T_4476 ? 16'h100 : _T_6313; // @[Mux.scala 31:69:@3263.4]
  assign _T_6315 = _T_4473 ? 16'h80 : _T_6314; // @[Mux.scala 31:69:@3264.4]
  assign _T_6316 = _T_4470 ? 16'h40 : _T_6315; // @[Mux.scala 31:69:@3265.4]
  assign _T_6317 = _T_4467 ? 16'h20 : _T_6316; // @[Mux.scala 31:69:@3266.4]
  assign _T_6318 = _T_4464 ? 16'h10 : _T_6317; // @[Mux.scala 31:69:@3267.4]
  assign _T_6319 = _T_4461 ? 16'h8 : _T_6318; // @[Mux.scala 31:69:@3268.4]
  assign _T_6320 = _T_4458 ? 16'h4 : _T_6319; // @[Mux.scala 31:69:@3269.4]
  assign _T_6321 = _T_4455 ? 16'h2 : _T_6320; // @[Mux.scala 31:69:@3270.4]
  assign _T_6322 = _T_4452 ? 16'h1 : _T_6321; // @[Mux.scala 31:69:@3271.4]
  assign _T_6323 = _T_6322[0]; // @[OneHot.scala 66:30:@3272.4]
  assign _T_6324 = _T_6322[1]; // @[OneHot.scala 66:30:@3273.4]
  assign _T_6325 = _T_6322[2]; // @[OneHot.scala 66:30:@3274.4]
  assign _T_6326 = _T_6322[3]; // @[OneHot.scala 66:30:@3275.4]
  assign _T_6327 = _T_6322[4]; // @[OneHot.scala 66:30:@3276.4]
  assign _T_6328 = _T_6322[5]; // @[OneHot.scala 66:30:@3277.4]
  assign _T_6329 = _T_6322[6]; // @[OneHot.scala 66:30:@3278.4]
  assign _T_6330 = _T_6322[7]; // @[OneHot.scala 66:30:@3279.4]
  assign _T_6331 = _T_6322[8]; // @[OneHot.scala 66:30:@3280.4]
  assign _T_6332 = _T_6322[9]; // @[OneHot.scala 66:30:@3281.4]
  assign _T_6333 = _T_6322[10]; // @[OneHot.scala 66:30:@3282.4]
  assign _T_6334 = _T_6322[11]; // @[OneHot.scala 66:30:@3283.4]
  assign _T_6335 = _T_6322[12]; // @[OneHot.scala 66:30:@3284.4]
  assign _T_6336 = _T_6322[13]; // @[OneHot.scala 66:30:@3285.4]
  assign _T_6337 = _T_6322[14]; // @[OneHot.scala 66:30:@3286.4]
  assign _T_6338 = _T_6322[15]; // @[OneHot.scala 66:30:@3287.4]
  assign _T_6379 = _T_4452 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3305.4]
  assign _T_6380 = _T_4449 ? 16'h4000 : _T_6379; // @[Mux.scala 31:69:@3306.4]
  assign _T_6381 = _T_4494 ? 16'h2000 : _T_6380; // @[Mux.scala 31:69:@3307.4]
  assign _T_6382 = _T_4491 ? 16'h1000 : _T_6381; // @[Mux.scala 31:69:@3308.4]
  assign _T_6383 = _T_4488 ? 16'h800 : _T_6382; // @[Mux.scala 31:69:@3309.4]
  assign _T_6384 = _T_4485 ? 16'h400 : _T_6383; // @[Mux.scala 31:69:@3310.4]
  assign _T_6385 = _T_4482 ? 16'h200 : _T_6384; // @[Mux.scala 31:69:@3311.4]
  assign _T_6386 = _T_4479 ? 16'h100 : _T_6385; // @[Mux.scala 31:69:@3312.4]
  assign _T_6387 = _T_4476 ? 16'h80 : _T_6386; // @[Mux.scala 31:69:@3313.4]
  assign _T_6388 = _T_4473 ? 16'h40 : _T_6387; // @[Mux.scala 31:69:@3314.4]
  assign _T_6389 = _T_4470 ? 16'h20 : _T_6388; // @[Mux.scala 31:69:@3315.4]
  assign _T_6390 = _T_4467 ? 16'h10 : _T_6389; // @[Mux.scala 31:69:@3316.4]
  assign _T_6391 = _T_4464 ? 16'h8 : _T_6390; // @[Mux.scala 31:69:@3317.4]
  assign _T_6392 = _T_4461 ? 16'h4 : _T_6391; // @[Mux.scala 31:69:@3318.4]
  assign _T_6393 = _T_4458 ? 16'h2 : _T_6392; // @[Mux.scala 31:69:@3319.4]
  assign _T_6394 = _T_4455 ? 16'h1 : _T_6393; // @[Mux.scala 31:69:@3320.4]
  assign _T_6395 = _T_6394[0]; // @[OneHot.scala 66:30:@3321.4]
  assign _T_6396 = _T_6394[1]; // @[OneHot.scala 66:30:@3322.4]
  assign _T_6397 = _T_6394[2]; // @[OneHot.scala 66:30:@3323.4]
  assign _T_6398 = _T_6394[3]; // @[OneHot.scala 66:30:@3324.4]
  assign _T_6399 = _T_6394[4]; // @[OneHot.scala 66:30:@3325.4]
  assign _T_6400 = _T_6394[5]; // @[OneHot.scala 66:30:@3326.4]
  assign _T_6401 = _T_6394[6]; // @[OneHot.scala 66:30:@3327.4]
  assign _T_6402 = _T_6394[7]; // @[OneHot.scala 66:30:@3328.4]
  assign _T_6403 = _T_6394[8]; // @[OneHot.scala 66:30:@3329.4]
  assign _T_6404 = _T_6394[9]; // @[OneHot.scala 66:30:@3330.4]
  assign _T_6405 = _T_6394[10]; // @[OneHot.scala 66:30:@3331.4]
  assign _T_6406 = _T_6394[11]; // @[OneHot.scala 66:30:@3332.4]
  assign _T_6407 = _T_6394[12]; // @[OneHot.scala 66:30:@3333.4]
  assign _T_6408 = _T_6394[13]; // @[OneHot.scala 66:30:@3334.4]
  assign _T_6409 = _T_6394[14]; // @[OneHot.scala 66:30:@3335.4]
  assign _T_6410 = _T_6394[15]; // @[OneHot.scala 66:30:@3336.4]
  assign _T_6451 = _T_4455 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3354.4]
  assign _T_6452 = _T_4452 ? 16'h4000 : _T_6451; // @[Mux.scala 31:69:@3355.4]
  assign _T_6453 = _T_4449 ? 16'h2000 : _T_6452; // @[Mux.scala 31:69:@3356.4]
  assign _T_6454 = _T_4494 ? 16'h1000 : _T_6453; // @[Mux.scala 31:69:@3357.4]
  assign _T_6455 = _T_4491 ? 16'h800 : _T_6454; // @[Mux.scala 31:69:@3358.4]
  assign _T_6456 = _T_4488 ? 16'h400 : _T_6455; // @[Mux.scala 31:69:@3359.4]
  assign _T_6457 = _T_4485 ? 16'h200 : _T_6456; // @[Mux.scala 31:69:@3360.4]
  assign _T_6458 = _T_4482 ? 16'h100 : _T_6457; // @[Mux.scala 31:69:@3361.4]
  assign _T_6459 = _T_4479 ? 16'h80 : _T_6458; // @[Mux.scala 31:69:@3362.4]
  assign _T_6460 = _T_4476 ? 16'h40 : _T_6459; // @[Mux.scala 31:69:@3363.4]
  assign _T_6461 = _T_4473 ? 16'h20 : _T_6460; // @[Mux.scala 31:69:@3364.4]
  assign _T_6462 = _T_4470 ? 16'h10 : _T_6461; // @[Mux.scala 31:69:@3365.4]
  assign _T_6463 = _T_4467 ? 16'h8 : _T_6462; // @[Mux.scala 31:69:@3366.4]
  assign _T_6464 = _T_4464 ? 16'h4 : _T_6463; // @[Mux.scala 31:69:@3367.4]
  assign _T_6465 = _T_4461 ? 16'h2 : _T_6464; // @[Mux.scala 31:69:@3368.4]
  assign _T_6466 = _T_4458 ? 16'h1 : _T_6465; // @[Mux.scala 31:69:@3369.4]
  assign _T_6467 = _T_6466[0]; // @[OneHot.scala 66:30:@3370.4]
  assign _T_6468 = _T_6466[1]; // @[OneHot.scala 66:30:@3371.4]
  assign _T_6469 = _T_6466[2]; // @[OneHot.scala 66:30:@3372.4]
  assign _T_6470 = _T_6466[3]; // @[OneHot.scala 66:30:@3373.4]
  assign _T_6471 = _T_6466[4]; // @[OneHot.scala 66:30:@3374.4]
  assign _T_6472 = _T_6466[5]; // @[OneHot.scala 66:30:@3375.4]
  assign _T_6473 = _T_6466[6]; // @[OneHot.scala 66:30:@3376.4]
  assign _T_6474 = _T_6466[7]; // @[OneHot.scala 66:30:@3377.4]
  assign _T_6475 = _T_6466[8]; // @[OneHot.scala 66:30:@3378.4]
  assign _T_6476 = _T_6466[9]; // @[OneHot.scala 66:30:@3379.4]
  assign _T_6477 = _T_6466[10]; // @[OneHot.scala 66:30:@3380.4]
  assign _T_6478 = _T_6466[11]; // @[OneHot.scala 66:30:@3381.4]
  assign _T_6479 = _T_6466[12]; // @[OneHot.scala 66:30:@3382.4]
  assign _T_6480 = _T_6466[13]; // @[OneHot.scala 66:30:@3383.4]
  assign _T_6481 = _T_6466[14]; // @[OneHot.scala 66:30:@3384.4]
  assign _T_6482 = _T_6466[15]; // @[OneHot.scala 66:30:@3385.4]
  assign _T_6523 = _T_4458 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3403.4]
  assign _T_6524 = _T_4455 ? 16'h4000 : _T_6523; // @[Mux.scala 31:69:@3404.4]
  assign _T_6525 = _T_4452 ? 16'h2000 : _T_6524; // @[Mux.scala 31:69:@3405.4]
  assign _T_6526 = _T_4449 ? 16'h1000 : _T_6525; // @[Mux.scala 31:69:@3406.4]
  assign _T_6527 = _T_4494 ? 16'h800 : _T_6526; // @[Mux.scala 31:69:@3407.4]
  assign _T_6528 = _T_4491 ? 16'h400 : _T_6527; // @[Mux.scala 31:69:@3408.4]
  assign _T_6529 = _T_4488 ? 16'h200 : _T_6528; // @[Mux.scala 31:69:@3409.4]
  assign _T_6530 = _T_4485 ? 16'h100 : _T_6529; // @[Mux.scala 31:69:@3410.4]
  assign _T_6531 = _T_4482 ? 16'h80 : _T_6530; // @[Mux.scala 31:69:@3411.4]
  assign _T_6532 = _T_4479 ? 16'h40 : _T_6531; // @[Mux.scala 31:69:@3412.4]
  assign _T_6533 = _T_4476 ? 16'h20 : _T_6532; // @[Mux.scala 31:69:@3413.4]
  assign _T_6534 = _T_4473 ? 16'h10 : _T_6533; // @[Mux.scala 31:69:@3414.4]
  assign _T_6535 = _T_4470 ? 16'h8 : _T_6534; // @[Mux.scala 31:69:@3415.4]
  assign _T_6536 = _T_4467 ? 16'h4 : _T_6535; // @[Mux.scala 31:69:@3416.4]
  assign _T_6537 = _T_4464 ? 16'h2 : _T_6536; // @[Mux.scala 31:69:@3417.4]
  assign _T_6538 = _T_4461 ? 16'h1 : _T_6537; // @[Mux.scala 31:69:@3418.4]
  assign _T_6539 = _T_6538[0]; // @[OneHot.scala 66:30:@3419.4]
  assign _T_6540 = _T_6538[1]; // @[OneHot.scala 66:30:@3420.4]
  assign _T_6541 = _T_6538[2]; // @[OneHot.scala 66:30:@3421.4]
  assign _T_6542 = _T_6538[3]; // @[OneHot.scala 66:30:@3422.4]
  assign _T_6543 = _T_6538[4]; // @[OneHot.scala 66:30:@3423.4]
  assign _T_6544 = _T_6538[5]; // @[OneHot.scala 66:30:@3424.4]
  assign _T_6545 = _T_6538[6]; // @[OneHot.scala 66:30:@3425.4]
  assign _T_6546 = _T_6538[7]; // @[OneHot.scala 66:30:@3426.4]
  assign _T_6547 = _T_6538[8]; // @[OneHot.scala 66:30:@3427.4]
  assign _T_6548 = _T_6538[9]; // @[OneHot.scala 66:30:@3428.4]
  assign _T_6549 = _T_6538[10]; // @[OneHot.scala 66:30:@3429.4]
  assign _T_6550 = _T_6538[11]; // @[OneHot.scala 66:30:@3430.4]
  assign _T_6551 = _T_6538[12]; // @[OneHot.scala 66:30:@3431.4]
  assign _T_6552 = _T_6538[13]; // @[OneHot.scala 66:30:@3432.4]
  assign _T_6553 = _T_6538[14]; // @[OneHot.scala 66:30:@3433.4]
  assign _T_6554 = _T_6538[15]; // @[OneHot.scala 66:30:@3434.4]
  assign _T_6595 = _T_4461 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3452.4]
  assign _T_6596 = _T_4458 ? 16'h4000 : _T_6595; // @[Mux.scala 31:69:@3453.4]
  assign _T_6597 = _T_4455 ? 16'h2000 : _T_6596; // @[Mux.scala 31:69:@3454.4]
  assign _T_6598 = _T_4452 ? 16'h1000 : _T_6597; // @[Mux.scala 31:69:@3455.4]
  assign _T_6599 = _T_4449 ? 16'h800 : _T_6598; // @[Mux.scala 31:69:@3456.4]
  assign _T_6600 = _T_4494 ? 16'h400 : _T_6599; // @[Mux.scala 31:69:@3457.4]
  assign _T_6601 = _T_4491 ? 16'h200 : _T_6600; // @[Mux.scala 31:69:@3458.4]
  assign _T_6602 = _T_4488 ? 16'h100 : _T_6601; // @[Mux.scala 31:69:@3459.4]
  assign _T_6603 = _T_4485 ? 16'h80 : _T_6602; // @[Mux.scala 31:69:@3460.4]
  assign _T_6604 = _T_4482 ? 16'h40 : _T_6603; // @[Mux.scala 31:69:@3461.4]
  assign _T_6605 = _T_4479 ? 16'h20 : _T_6604; // @[Mux.scala 31:69:@3462.4]
  assign _T_6606 = _T_4476 ? 16'h10 : _T_6605; // @[Mux.scala 31:69:@3463.4]
  assign _T_6607 = _T_4473 ? 16'h8 : _T_6606; // @[Mux.scala 31:69:@3464.4]
  assign _T_6608 = _T_4470 ? 16'h4 : _T_6607; // @[Mux.scala 31:69:@3465.4]
  assign _T_6609 = _T_4467 ? 16'h2 : _T_6608; // @[Mux.scala 31:69:@3466.4]
  assign _T_6610 = _T_4464 ? 16'h1 : _T_6609; // @[Mux.scala 31:69:@3467.4]
  assign _T_6611 = _T_6610[0]; // @[OneHot.scala 66:30:@3468.4]
  assign _T_6612 = _T_6610[1]; // @[OneHot.scala 66:30:@3469.4]
  assign _T_6613 = _T_6610[2]; // @[OneHot.scala 66:30:@3470.4]
  assign _T_6614 = _T_6610[3]; // @[OneHot.scala 66:30:@3471.4]
  assign _T_6615 = _T_6610[4]; // @[OneHot.scala 66:30:@3472.4]
  assign _T_6616 = _T_6610[5]; // @[OneHot.scala 66:30:@3473.4]
  assign _T_6617 = _T_6610[6]; // @[OneHot.scala 66:30:@3474.4]
  assign _T_6618 = _T_6610[7]; // @[OneHot.scala 66:30:@3475.4]
  assign _T_6619 = _T_6610[8]; // @[OneHot.scala 66:30:@3476.4]
  assign _T_6620 = _T_6610[9]; // @[OneHot.scala 66:30:@3477.4]
  assign _T_6621 = _T_6610[10]; // @[OneHot.scala 66:30:@3478.4]
  assign _T_6622 = _T_6610[11]; // @[OneHot.scala 66:30:@3479.4]
  assign _T_6623 = _T_6610[12]; // @[OneHot.scala 66:30:@3480.4]
  assign _T_6624 = _T_6610[13]; // @[OneHot.scala 66:30:@3481.4]
  assign _T_6625 = _T_6610[14]; // @[OneHot.scala 66:30:@3482.4]
  assign _T_6626 = _T_6610[15]; // @[OneHot.scala 66:30:@3483.4]
  assign _T_6667 = _T_4464 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3501.4]
  assign _T_6668 = _T_4461 ? 16'h4000 : _T_6667; // @[Mux.scala 31:69:@3502.4]
  assign _T_6669 = _T_4458 ? 16'h2000 : _T_6668; // @[Mux.scala 31:69:@3503.4]
  assign _T_6670 = _T_4455 ? 16'h1000 : _T_6669; // @[Mux.scala 31:69:@3504.4]
  assign _T_6671 = _T_4452 ? 16'h800 : _T_6670; // @[Mux.scala 31:69:@3505.4]
  assign _T_6672 = _T_4449 ? 16'h400 : _T_6671; // @[Mux.scala 31:69:@3506.4]
  assign _T_6673 = _T_4494 ? 16'h200 : _T_6672; // @[Mux.scala 31:69:@3507.4]
  assign _T_6674 = _T_4491 ? 16'h100 : _T_6673; // @[Mux.scala 31:69:@3508.4]
  assign _T_6675 = _T_4488 ? 16'h80 : _T_6674; // @[Mux.scala 31:69:@3509.4]
  assign _T_6676 = _T_4485 ? 16'h40 : _T_6675; // @[Mux.scala 31:69:@3510.4]
  assign _T_6677 = _T_4482 ? 16'h20 : _T_6676; // @[Mux.scala 31:69:@3511.4]
  assign _T_6678 = _T_4479 ? 16'h10 : _T_6677; // @[Mux.scala 31:69:@3512.4]
  assign _T_6679 = _T_4476 ? 16'h8 : _T_6678; // @[Mux.scala 31:69:@3513.4]
  assign _T_6680 = _T_4473 ? 16'h4 : _T_6679; // @[Mux.scala 31:69:@3514.4]
  assign _T_6681 = _T_4470 ? 16'h2 : _T_6680; // @[Mux.scala 31:69:@3515.4]
  assign _T_6682 = _T_4467 ? 16'h1 : _T_6681; // @[Mux.scala 31:69:@3516.4]
  assign _T_6683 = _T_6682[0]; // @[OneHot.scala 66:30:@3517.4]
  assign _T_6684 = _T_6682[1]; // @[OneHot.scala 66:30:@3518.4]
  assign _T_6685 = _T_6682[2]; // @[OneHot.scala 66:30:@3519.4]
  assign _T_6686 = _T_6682[3]; // @[OneHot.scala 66:30:@3520.4]
  assign _T_6687 = _T_6682[4]; // @[OneHot.scala 66:30:@3521.4]
  assign _T_6688 = _T_6682[5]; // @[OneHot.scala 66:30:@3522.4]
  assign _T_6689 = _T_6682[6]; // @[OneHot.scala 66:30:@3523.4]
  assign _T_6690 = _T_6682[7]; // @[OneHot.scala 66:30:@3524.4]
  assign _T_6691 = _T_6682[8]; // @[OneHot.scala 66:30:@3525.4]
  assign _T_6692 = _T_6682[9]; // @[OneHot.scala 66:30:@3526.4]
  assign _T_6693 = _T_6682[10]; // @[OneHot.scala 66:30:@3527.4]
  assign _T_6694 = _T_6682[11]; // @[OneHot.scala 66:30:@3528.4]
  assign _T_6695 = _T_6682[12]; // @[OneHot.scala 66:30:@3529.4]
  assign _T_6696 = _T_6682[13]; // @[OneHot.scala 66:30:@3530.4]
  assign _T_6697 = _T_6682[14]; // @[OneHot.scala 66:30:@3531.4]
  assign _T_6698 = _T_6682[15]; // @[OneHot.scala 66:30:@3532.4]
  assign _T_6739 = _T_4467 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3550.4]
  assign _T_6740 = _T_4464 ? 16'h4000 : _T_6739; // @[Mux.scala 31:69:@3551.4]
  assign _T_6741 = _T_4461 ? 16'h2000 : _T_6740; // @[Mux.scala 31:69:@3552.4]
  assign _T_6742 = _T_4458 ? 16'h1000 : _T_6741; // @[Mux.scala 31:69:@3553.4]
  assign _T_6743 = _T_4455 ? 16'h800 : _T_6742; // @[Mux.scala 31:69:@3554.4]
  assign _T_6744 = _T_4452 ? 16'h400 : _T_6743; // @[Mux.scala 31:69:@3555.4]
  assign _T_6745 = _T_4449 ? 16'h200 : _T_6744; // @[Mux.scala 31:69:@3556.4]
  assign _T_6746 = _T_4494 ? 16'h100 : _T_6745; // @[Mux.scala 31:69:@3557.4]
  assign _T_6747 = _T_4491 ? 16'h80 : _T_6746; // @[Mux.scala 31:69:@3558.4]
  assign _T_6748 = _T_4488 ? 16'h40 : _T_6747; // @[Mux.scala 31:69:@3559.4]
  assign _T_6749 = _T_4485 ? 16'h20 : _T_6748; // @[Mux.scala 31:69:@3560.4]
  assign _T_6750 = _T_4482 ? 16'h10 : _T_6749; // @[Mux.scala 31:69:@3561.4]
  assign _T_6751 = _T_4479 ? 16'h8 : _T_6750; // @[Mux.scala 31:69:@3562.4]
  assign _T_6752 = _T_4476 ? 16'h4 : _T_6751; // @[Mux.scala 31:69:@3563.4]
  assign _T_6753 = _T_4473 ? 16'h2 : _T_6752; // @[Mux.scala 31:69:@3564.4]
  assign _T_6754 = _T_4470 ? 16'h1 : _T_6753; // @[Mux.scala 31:69:@3565.4]
  assign _T_6755 = _T_6754[0]; // @[OneHot.scala 66:30:@3566.4]
  assign _T_6756 = _T_6754[1]; // @[OneHot.scala 66:30:@3567.4]
  assign _T_6757 = _T_6754[2]; // @[OneHot.scala 66:30:@3568.4]
  assign _T_6758 = _T_6754[3]; // @[OneHot.scala 66:30:@3569.4]
  assign _T_6759 = _T_6754[4]; // @[OneHot.scala 66:30:@3570.4]
  assign _T_6760 = _T_6754[5]; // @[OneHot.scala 66:30:@3571.4]
  assign _T_6761 = _T_6754[6]; // @[OneHot.scala 66:30:@3572.4]
  assign _T_6762 = _T_6754[7]; // @[OneHot.scala 66:30:@3573.4]
  assign _T_6763 = _T_6754[8]; // @[OneHot.scala 66:30:@3574.4]
  assign _T_6764 = _T_6754[9]; // @[OneHot.scala 66:30:@3575.4]
  assign _T_6765 = _T_6754[10]; // @[OneHot.scala 66:30:@3576.4]
  assign _T_6766 = _T_6754[11]; // @[OneHot.scala 66:30:@3577.4]
  assign _T_6767 = _T_6754[12]; // @[OneHot.scala 66:30:@3578.4]
  assign _T_6768 = _T_6754[13]; // @[OneHot.scala 66:30:@3579.4]
  assign _T_6769 = _T_6754[14]; // @[OneHot.scala 66:30:@3580.4]
  assign _T_6770 = _T_6754[15]; // @[OneHot.scala 66:30:@3581.4]
  assign _T_6811 = _T_4470 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3599.4]
  assign _T_6812 = _T_4467 ? 16'h4000 : _T_6811; // @[Mux.scala 31:69:@3600.4]
  assign _T_6813 = _T_4464 ? 16'h2000 : _T_6812; // @[Mux.scala 31:69:@3601.4]
  assign _T_6814 = _T_4461 ? 16'h1000 : _T_6813; // @[Mux.scala 31:69:@3602.4]
  assign _T_6815 = _T_4458 ? 16'h800 : _T_6814; // @[Mux.scala 31:69:@3603.4]
  assign _T_6816 = _T_4455 ? 16'h400 : _T_6815; // @[Mux.scala 31:69:@3604.4]
  assign _T_6817 = _T_4452 ? 16'h200 : _T_6816; // @[Mux.scala 31:69:@3605.4]
  assign _T_6818 = _T_4449 ? 16'h100 : _T_6817; // @[Mux.scala 31:69:@3606.4]
  assign _T_6819 = _T_4494 ? 16'h80 : _T_6818; // @[Mux.scala 31:69:@3607.4]
  assign _T_6820 = _T_4491 ? 16'h40 : _T_6819; // @[Mux.scala 31:69:@3608.4]
  assign _T_6821 = _T_4488 ? 16'h20 : _T_6820; // @[Mux.scala 31:69:@3609.4]
  assign _T_6822 = _T_4485 ? 16'h10 : _T_6821; // @[Mux.scala 31:69:@3610.4]
  assign _T_6823 = _T_4482 ? 16'h8 : _T_6822; // @[Mux.scala 31:69:@3611.4]
  assign _T_6824 = _T_4479 ? 16'h4 : _T_6823; // @[Mux.scala 31:69:@3612.4]
  assign _T_6825 = _T_4476 ? 16'h2 : _T_6824; // @[Mux.scala 31:69:@3613.4]
  assign _T_6826 = _T_4473 ? 16'h1 : _T_6825; // @[Mux.scala 31:69:@3614.4]
  assign _T_6827 = _T_6826[0]; // @[OneHot.scala 66:30:@3615.4]
  assign _T_6828 = _T_6826[1]; // @[OneHot.scala 66:30:@3616.4]
  assign _T_6829 = _T_6826[2]; // @[OneHot.scala 66:30:@3617.4]
  assign _T_6830 = _T_6826[3]; // @[OneHot.scala 66:30:@3618.4]
  assign _T_6831 = _T_6826[4]; // @[OneHot.scala 66:30:@3619.4]
  assign _T_6832 = _T_6826[5]; // @[OneHot.scala 66:30:@3620.4]
  assign _T_6833 = _T_6826[6]; // @[OneHot.scala 66:30:@3621.4]
  assign _T_6834 = _T_6826[7]; // @[OneHot.scala 66:30:@3622.4]
  assign _T_6835 = _T_6826[8]; // @[OneHot.scala 66:30:@3623.4]
  assign _T_6836 = _T_6826[9]; // @[OneHot.scala 66:30:@3624.4]
  assign _T_6837 = _T_6826[10]; // @[OneHot.scala 66:30:@3625.4]
  assign _T_6838 = _T_6826[11]; // @[OneHot.scala 66:30:@3626.4]
  assign _T_6839 = _T_6826[12]; // @[OneHot.scala 66:30:@3627.4]
  assign _T_6840 = _T_6826[13]; // @[OneHot.scala 66:30:@3628.4]
  assign _T_6841 = _T_6826[14]; // @[OneHot.scala 66:30:@3629.4]
  assign _T_6842 = _T_6826[15]; // @[OneHot.scala 66:30:@3630.4]
  assign _T_6883 = _T_4473 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3648.4]
  assign _T_6884 = _T_4470 ? 16'h4000 : _T_6883; // @[Mux.scala 31:69:@3649.4]
  assign _T_6885 = _T_4467 ? 16'h2000 : _T_6884; // @[Mux.scala 31:69:@3650.4]
  assign _T_6886 = _T_4464 ? 16'h1000 : _T_6885; // @[Mux.scala 31:69:@3651.4]
  assign _T_6887 = _T_4461 ? 16'h800 : _T_6886; // @[Mux.scala 31:69:@3652.4]
  assign _T_6888 = _T_4458 ? 16'h400 : _T_6887; // @[Mux.scala 31:69:@3653.4]
  assign _T_6889 = _T_4455 ? 16'h200 : _T_6888; // @[Mux.scala 31:69:@3654.4]
  assign _T_6890 = _T_4452 ? 16'h100 : _T_6889; // @[Mux.scala 31:69:@3655.4]
  assign _T_6891 = _T_4449 ? 16'h80 : _T_6890; // @[Mux.scala 31:69:@3656.4]
  assign _T_6892 = _T_4494 ? 16'h40 : _T_6891; // @[Mux.scala 31:69:@3657.4]
  assign _T_6893 = _T_4491 ? 16'h20 : _T_6892; // @[Mux.scala 31:69:@3658.4]
  assign _T_6894 = _T_4488 ? 16'h10 : _T_6893; // @[Mux.scala 31:69:@3659.4]
  assign _T_6895 = _T_4485 ? 16'h8 : _T_6894; // @[Mux.scala 31:69:@3660.4]
  assign _T_6896 = _T_4482 ? 16'h4 : _T_6895; // @[Mux.scala 31:69:@3661.4]
  assign _T_6897 = _T_4479 ? 16'h2 : _T_6896; // @[Mux.scala 31:69:@3662.4]
  assign _T_6898 = _T_4476 ? 16'h1 : _T_6897; // @[Mux.scala 31:69:@3663.4]
  assign _T_6899 = _T_6898[0]; // @[OneHot.scala 66:30:@3664.4]
  assign _T_6900 = _T_6898[1]; // @[OneHot.scala 66:30:@3665.4]
  assign _T_6901 = _T_6898[2]; // @[OneHot.scala 66:30:@3666.4]
  assign _T_6902 = _T_6898[3]; // @[OneHot.scala 66:30:@3667.4]
  assign _T_6903 = _T_6898[4]; // @[OneHot.scala 66:30:@3668.4]
  assign _T_6904 = _T_6898[5]; // @[OneHot.scala 66:30:@3669.4]
  assign _T_6905 = _T_6898[6]; // @[OneHot.scala 66:30:@3670.4]
  assign _T_6906 = _T_6898[7]; // @[OneHot.scala 66:30:@3671.4]
  assign _T_6907 = _T_6898[8]; // @[OneHot.scala 66:30:@3672.4]
  assign _T_6908 = _T_6898[9]; // @[OneHot.scala 66:30:@3673.4]
  assign _T_6909 = _T_6898[10]; // @[OneHot.scala 66:30:@3674.4]
  assign _T_6910 = _T_6898[11]; // @[OneHot.scala 66:30:@3675.4]
  assign _T_6911 = _T_6898[12]; // @[OneHot.scala 66:30:@3676.4]
  assign _T_6912 = _T_6898[13]; // @[OneHot.scala 66:30:@3677.4]
  assign _T_6913 = _T_6898[14]; // @[OneHot.scala 66:30:@3678.4]
  assign _T_6914 = _T_6898[15]; // @[OneHot.scala 66:30:@3679.4]
  assign _T_6955 = _T_4476 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3697.4]
  assign _T_6956 = _T_4473 ? 16'h4000 : _T_6955; // @[Mux.scala 31:69:@3698.4]
  assign _T_6957 = _T_4470 ? 16'h2000 : _T_6956; // @[Mux.scala 31:69:@3699.4]
  assign _T_6958 = _T_4467 ? 16'h1000 : _T_6957; // @[Mux.scala 31:69:@3700.4]
  assign _T_6959 = _T_4464 ? 16'h800 : _T_6958; // @[Mux.scala 31:69:@3701.4]
  assign _T_6960 = _T_4461 ? 16'h400 : _T_6959; // @[Mux.scala 31:69:@3702.4]
  assign _T_6961 = _T_4458 ? 16'h200 : _T_6960; // @[Mux.scala 31:69:@3703.4]
  assign _T_6962 = _T_4455 ? 16'h100 : _T_6961; // @[Mux.scala 31:69:@3704.4]
  assign _T_6963 = _T_4452 ? 16'h80 : _T_6962; // @[Mux.scala 31:69:@3705.4]
  assign _T_6964 = _T_4449 ? 16'h40 : _T_6963; // @[Mux.scala 31:69:@3706.4]
  assign _T_6965 = _T_4494 ? 16'h20 : _T_6964; // @[Mux.scala 31:69:@3707.4]
  assign _T_6966 = _T_4491 ? 16'h10 : _T_6965; // @[Mux.scala 31:69:@3708.4]
  assign _T_6967 = _T_4488 ? 16'h8 : _T_6966; // @[Mux.scala 31:69:@3709.4]
  assign _T_6968 = _T_4485 ? 16'h4 : _T_6967; // @[Mux.scala 31:69:@3710.4]
  assign _T_6969 = _T_4482 ? 16'h2 : _T_6968; // @[Mux.scala 31:69:@3711.4]
  assign _T_6970 = _T_4479 ? 16'h1 : _T_6969; // @[Mux.scala 31:69:@3712.4]
  assign _T_6971 = _T_6970[0]; // @[OneHot.scala 66:30:@3713.4]
  assign _T_6972 = _T_6970[1]; // @[OneHot.scala 66:30:@3714.4]
  assign _T_6973 = _T_6970[2]; // @[OneHot.scala 66:30:@3715.4]
  assign _T_6974 = _T_6970[3]; // @[OneHot.scala 66:30:@3716.4]
  assign _T_6975 = _T_6970[4]; // @[OneHot.scala 66:30:@3717.4]
  assign _T_6976 = _T_6970[5]; // @[OneHot.scala 66:30:@3718.4]
  assign _T_6977 = _T_6970[6]; // @[OneHot.scala 66:30:@3719.4]
  assign _T_6978 = _T_6970[7]; // @[OneHot.scala 66:30:@3720.4]
  assign _T_6979 = _T_6970[8]; // @[OneHot.scala 66:30:@3721.4]
  assign _T_6980 = _T_6970[9]; // @[OneHot.scala 66:30:@3722.4]
  assign _T_6981 = _T_6970[10]; // @[OneHot.scala 66:30:@3723.4]
  assign _T_6982 = _T_6970[11]; // @[OneHot.scala 66:30:@3724.4]
  assign _T_6983 = _T_6970[12]; // @[OneHot.scala 66:30:@3725.4]
  assign _T_6984 = _T_6970[13]; // @[OneHot.scala 66:30:@3726.4]
  assign _T_6985 = _T_6970[14]; // @[OneHot.scala 66:30:@3727.4]
  assign _T_6986 = _T_6970[15]; // @[OneHot.scala 66:30:@3728.4]
  assign _T_7027 = _T_4479 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3746.4]
  assign _T_7028 = _T_4476 ? 16'h4000 : _T_7027; // @[Mux.scala 31:69:@3747.4]
  assign _T_7029 = _T_4473 ? 16'h2000 : _T_7028; // @[Mux.scala 31:69:@3748.4]
  assign _T_7030 = _T_4470 ? 16'h1000 : _T_7029; // @[Mux.scala 31:69:@3749.4]
  assign _T_7031 = _T_4467 ? 16'h800 : _T_7030; // @[Mux.scala 31:69:@3750.4]
  assign _T_7032 = _T_4464 ? 16'h400 : _T_7031; // @[Mux.scala 31:69:@3751.4]
  assign _T_7033 = _T_4461 ? 16'h200 : _T_7032; // @[Mux.scala 31:69:@3752.4]
  assign _T_7034 = _T_4458 ? 16'h100 : _T_7033; // @[Mux.scala 31:69:@3753.4]
  assign _T_7035 = _T_4455 ? 16'h80 : _T_7034; // @[Mux.scala 31:69:@3754.4]
  assign _T_7036 = _T_4452 ? 16'h40 : _T_7035; // @[Mux.scala 31:69:@3755.4]
  assign _T_7037 = _T_4449 ? 16'h20 : _T_7036; // @[Mux.scala 31:69:@3756.4]
  assign _T_7038 = _T_4494 ? 16'h10 : _T_7037; // @[Mux.scala 31:69:@3757.4]
  assign _T_7039 = _T_4491 ? 16'h8 : _T_7038; // @[Mux.scala 31:69:@3758.4]
  assign _T_7040 = _T_4488 ? 16'h4 : _T_7039; // @[Mux.scala 31:69:@3759.4]
  assign _T_7041 = _T_4485 ? 16'h2 : _T_7040; // @[Mux.scala 31:69:@3760.4]
  assign _T_7042 = _T_4482 ? 16'h1 : _T_7041; // @[Mux.scala 31:69:@3761.4]
  assign _T_7043 = _T_7042[0]; // @[OneHot.scala 66:30:@3762.4]
  assign _T_7044 = _T_7042[1]; // @[OneHot.scala 66:30:@3763.4]
  assign _T_7045 = _T_7042[2]; // @[OneHot.scala 66:30:@3764.4]
  assign _T_7046 = _T_7042[3]; // @[OneHot.scala 66:30:@3765.4]
  assign _T_7047 = _T_7042[4]; // @[OneHot.scala 66:30:@3766.4]
  assign _T_7048 = _T_7042[5]; // @[OneHot.scala 66:30:@3767.4]
  assign _T_7049 = _T_7042[6]; // @[OneHot.scala 66:30:@3768.4]
  assign _T_7050 = _T_7042[7]; // @[OneHot.scala 66:30:@3769.4]
  assign _T_7051 = _T_7042[8]; // @[OneHot.scala 66:30:@3770.4]
  assign _T_7052 = _T_7042[9]; // @[OneHot.scala 66:30:@3771.4]
  assign _T_7053 = _T_7042[10]; // @[OneHot.scala 66:30:@3772.4]
  assign _T_7054 = _T_7042[11]; // @[OneHot.scala 66:30:@3773.4]
  assign _T_7055 = _T_7042[12]; // @[OneHot.scala 66:30:@3774.4]
  assign _T_7056 = _T_7042[13]; // @[OneHot.scala 66:30:@3775.4]
  assign _T_7057 = _T_7042[14]; // @[OneHot.scala 66:30:@3776.4]
  assign _T_7058 = _T_7042[15]; // @[OneHot.scala 66:30:@3777.4]
  assign _T_7099 = _T_4482 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3795.4]
  assign _T_7100 = _T_4479 ? 16'h4000 : _T_7099; // @[Mux.scala 31:69:@3796.4]
  assign _T_7101 = _T_4476 ? 16'h2000 : _T_7100; // @[Mux.scala 31:69:@3797.4]
  assign _T_7102 = _T_4473 ? 16'h1000 : _T_7101; // @[Mux.scala 31:69:@3798.4]
  assign _T_7103 = _T_4470 ? 16'h800 : _T_7102; // @[Mux.scala 31:69:@3799.4]
  assign _T_7104 = _T_4467 ? 16'h400 : _T_7103; // @[Mux.scala 31:69:@3800.4]
  assign _T_7105 = _T_4464 ? 16'h200 : _T_7104; // @[Mux.scala 31:69:@3801.4]
  assign _T_7106 = _T_4461 ? 16'h100 : _T_7105; // @[Mux.scala 31:69:@3802.4]
  assign _T_7107 = _T_4458 ? 16'h80 : _T_7106; // @[Mux.scala 31:69:@3803.4]
  assign _T_7108 = _T_4455 ? 16'h40 : _T_7107; // @[Mux.scala 31:69:@3804.4]
  assign _T_7109 = _T_4452 ? 16'h20 : _T_7108; // @[Mux.scala 31:69:@3805.4]
  assign _T_7110 = _T_4449 ? 16'h10 : _T_7109; // @[Mux.scala 31:69:@3806.4]
  assign _T_7111 = _T_4494 ? 16'h8 : _T_7110; // @[Mux.scala 31:69:@3807.4]
  assign _T_7112 = _T_4491 ? 16'h4 : _T_7111; // @[Mux.scala 31:69:@3808.4]
  assign _T_7113 = _T_4488 ? 16'h2 : _T_7112; // @[Mux.scala 31:69:@3809.4]
  assign _T_7114 = _T_4485 ? 16'h1 : _T_7113; // @[Mux.scala 31:69:@3810.4]
  assign _T_7115 = _T_7114[0]; // @[OneHot.scala 66:30:@3811.4]
  assign _T_7116 = _T_7114[1]; // @[OneHot.scala 66:30:@3812.4]
  assign _T_7117 = _T_7114[2]; // @[OneHot.scala 66:30:@3813.4]
  assign _T_7118 = _T_7114[3]; // @[OneHot.scala 66:30:@3814.4]
  assign _T_7119 = _T_7114[4]; // @[OneHot.scala 66:30:@3815.4]
  assign _T_7120 = _T_7114[5]; // @[OneHot.scala 66:30:@3816.4]
  assign _T_7121 = _T_7114[6]; // @[OneHot.scala 66:30:@3817.4]
  assign _T_7122 = _T_7114[7]; // @[OneHot.scala 66:30:@3818.4]
  assign _T_7123 = _T_7114[8]; // @[OneHot.scala 66:30:@3819.4]
  assign _T_7124 = _T_7114[9]; // @[OneHot.scala 66:30:@3820.4]
  assign _T_7125 = _T_7114[10]; // @[OneHot.scala 66:30:@3821.4]
  assign _T_7126 = _T_7114[11]; // @[OneHot.scala 66:30:@3822.4]
  assign _T_7127 = _T_7114[12]; // @[OneHot.scala 66:30:@3823.4]
  assign _T_7128 = _T_7114[13]; // @[OneHot.scala 66:30:@3824.4]
  assign _T_7129 = _T_7114[14]; // @[OneHot.scala 66:30:@3825.4]
  assign _T_7130 = _T_7114[15]; // @[OneHot.scala 66:30:@3826.4]
  assign _T_7171 = _T_4485 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3844.4]
  assign _T_7172 = _T_4482 ? 16'h4000 : _T_7171; // @[Mux.scala 31:69:@3845.4]
  assign _T_7173 = _T_4479 ? 16'h2000 : _T_7172; // @[Mux.scala 31:69:@3846.4]
  assign _T_7174 = _T_4476 ? 16'h1000 : _T_7173; // @[Mux.scala 31:69:@3847.4]
  assign _T_7175 = _T_4473 ? 16'h800 : _T_7174; // @[Mux.scala 31:69:@3848.4]
  assign _T_7176 = _T_4470 ? 16'h400 : _T_7175; // @[Mux.scala 31:69:@3849.4]
  assign _T_7177 = _T_4467 ? 16'h200 : _T_7176; // @[Mux.scala 31:69:@3850.4]
  assign _T_7178 = _T_4464 ? 16'h100 : _T_7177; // @[Mux.scala 31:69:@3851.4]
  assign _T_7179 = _T_4461 ? 16'h80 : _T_7178; // @[Mux.scala 31:69:@3852.4]
  assign _T_7180 = _T_4458 ? 16'h40 : _T_7179; // @[Mux.scala 31:69:@3853.4]
  assign _T_7181 = _T_4455 ? 16'h20 : _T_7180; // @[Mux.scala 31:69:@3854.4]
  assign _T_7182 = _T_4452 ? 16'h10 : _T_7181; // @[Mux.scala 31:69:@3855.4]
  assign _T_7183 = _T_4449 ? 16'h8 : _T_7182; // @[Mux.scala 31:69:@3856.4]
  assign _T_7184 = _T_4494 ? 16'h4 : _T_7183; // @[Mux.scala 31:69:@3857.4]
  assign _T_7185 = _T_4491 ? 16'h2 : _T_7184; // @[Mux.scala 31:69:@3858.4]
  assign _T_7186 = _T_4488 ? 16'h1 : _T_7185; // @[Mux.scala 31:69:@3859.4]
  assign _T_7187 = _T_7186[0]; // @[OneHot.scala 66:30:@3860.4]
  assign _T_7188 = _T_7186[1]; // @[OneHot.scala 66:30:@3861.4]
  assign _T_7189 = _T_7186[2]; // @[OneHot.scala 66:30:@3862.4]
  assign _T_7190 = _T_7186[3]; // @[OneHot.scala 66:30:@3863.4]
  assign _T_7191 = _T_7186[4]; // @[OneHot.scala 66:30:@3864.4]
  assign _T_7192 = _T_7186[5]; // @[OneHot.scala 66:30:@3865.4]
  assign _T_7193 = _T_7186[6]; // @[OneHot.scala 66:30:@3866.4]
  assign _T_7194 = _T_7186[7]; // @[OneHot.scala 66:30:@3867.4]
  assign _T_7195 = _T_7186[8]; // @[OneHot.scala 66:30:@3868.4]
  assign _T_7196 = _T_7186[9]; // @[OneHot.scala 66:30:@3869.4]
  assign _T_7197 = _T_7186[10]; // @[OneHot.scala 66:30:@3870.4]
  assign _T_7198 = _T_7186[11]; // @[OneHot.scala 66:30:@3871.4]
  assign _T_7199 = _T_7186[12]; // @[OneHot.scala 66:30:@3872.4]
  assign _T_7200 = _T_7186[13]; // @[OneHot.scala 66:30:@3873.4]
  assign _T_7201 = _T_7186[14]; // @[OneHot.scala 66:30:@3874.4]
  assign _T_7202 = _T_7186[15]; // @[OneHot.scala 66:30:@3875.4]
  assign _T_7243 = _T_4488 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3893.4]
  assign _T_7244 = _T_4485 ? 16'h4000 : _T_7243; // @[Mux.scala 31:69:@3894.4]
  assign _T_7245 = _T_4482 ? 16'h2000 : _T_7244; // @[Mux.scala 31:69:@3895.4]
  assign _T_7246 = _T_4479 ? 16'h1000 : _T_7245; // @[Mux.scala 31:69:@3896.4]
  assign _T_7247 = _T_4476 ? 16'h800 : _T_7246; // @[Mux.scala 31:69:@3897.4]
  assign _T_7248 = _T_4473 ? 16'h400 : _T_7247; // @[Mux.scala 31:69:@3898.4]
  assign _T_7249 = _T_4470 ? 16'h200 : _T_7248; // @[Mux.scala 31:69:@3899.4]
  assign _T_7250 = _T_4467 ? 16'h100 : _T_7249; // @[Mux.scala 31:69:@3900.4]
  assign _T_7251 = _T_4464 ? 16'h80 : _T_7250; // @[Mux.scala 31:69:@3901.4]
  assign _T_7252 = _T_4461 ? 16'h40 : _T_7251; // @[Mux.scala 31:69:@3902.4]
  assign _T_7253 = _T_4458 ? 16'h20 : _T_7252; // @[Mux.scala 31:69:@3903.4]
  assign _T_7254 = _T_4455 ? 16'h10 : _T_7253; // @[Mux.scala 31:69:@3904.4]
  assign _T_7255 = _T_4452 ? 16'h8 : _T_7254; // @[Mux.scala 31:69:@3905.4]
  assign _T_7256 = _T_4449 ? 16'h4 : _T_7255; // @[Mux.scala 31:69:@3906.4]
  assign _T_7257 = _T_4494 ? 16'h2 : _T_7256; // @[Mux.scala 31:69:@3907.4]
  assign _T_7258 = _T_4491 ? 16'h1 : _T_7257; // @[Mux.scala 31:69:@3908.4]
  assign _T_7259 = _T_7258[0]; // @[OneHot.scala 66:30:@3909.4]
  assign _T_7260 = _T_7258[1]; // @[OneHot.scala 66:30:@3910.4]
  assign _T_7261 = _T_7258[2]; // @[OneHot.scala 66:30:@3911.4]
  assign _T_7262 = _T_7258[3]; // @[OneHot.scala 66:30:@3912.4]
  assign _T_7263 = _T_7258[4]; // @[OneHot.scala 66:30:@3913.4]
  assign _T_7264 = _T_7258[5]; // @[OneHot.scala 66:30:@3914.4]
  assign _T_7265 = _T_7258[6]; // @[OneHot.scala 66:30:@3915.4]
  assign _T_7266 = _T_7258[7]; // @[OneHot.scala 66:30:@3916.4]
  assign _T_7267 = _T_7258[8]; // @[OneHot.scala 66:30:@3917.4]
  assign _T_7268 = _T_7258[9]; // @[OneHot.scala 66:30:@3918.4]
  assign _T_7269 = _T_7258[10]; // @[OneHot.scala 66:30:@3919.4]
  assign _T_7270 = _T_7258[11]; // @[OneHot.scala 66:30:@3920.4]
  assign _T_7271 = _T_7258[12]; // @[OneHot.scala 66:30:@3921.4]
  assign _T_7272 = _T_7258[13]; // @[OneHot.scala 66:30:@3922.4]
  assign _T_7273 = _T_7258[14]; // @[OneHot.scala 66:30:@3923.4]
  assign _T_7274 = _T_7258[15]; // @[OneHot.scala 66:30:@3924.4]
  assign _T_7315 = _T_4491 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3942.4]
  assign _T_7316 = _T_4488 ? 16'h4000 : _T_7315; // @[Mux.scala 31:69:@3943.4]
  assign _T_7317 = _T_4485 ? 16'h2000 : _T_7316; // @[Mux.scala 31:69:@3944.4]
  assign _T_7318 = _T_4482 ? 16'h1000 : _T_7317; // @[Mux.scala 31:69:@3945.4]
  assign _T_7319 = _T_4479 ? 16'h800 : _T_7318; // @[Mux.scala 31:69:@3946.4]
  assign _T_7320 = _T_4476 ? 16'h400 : _T_7319; // @[Mux.scala 31:69:@3947.4]
  assign _T_7321 = _T_4473 ? 16'h200 : _T_7320; // @[Mux.scala 31:69:@3948.4]
  assign _T_7322 = _T_4470 ? 16'h100 : _T_7321; // @[Mux.scala 31:69:@3949.4]
  assign _T_7323 = _T_4467 ? 16'h80 : _T_7322; // @[Mux.scala 31:69:@3950.4]
  assign _T_7324 = _T_4464 ? 16'h40 : _T_7323; // @[Mux.scala 31:69:@3951.4]
  assign _T_7325 = _T_4461 ? 16'h20 : _T_7324; // @[Mux.scala 31:69:@3952.4]
  assign _T_7326 = _T_4458 ? 16'h10 : _T_7325; // @[Mux.scala 31:69:@3953.4]
  assign _T_7327 = _T_4455 ? 16'h8 : _T_7326; // @[Mux.scala 31:69:@3954.4]
  assign _T_7328 = _T_4452 ? 16'h4 : _T_7327; // @[Mux.scala 31:69:@3955.4]
  assign _T_7329 = _T_4449 ? 16'h2 : _T_7328; // @[Mux.scala 31:69:@3956.4]
  assign _T_7330 = _T_4494 ? 16'h1 : _T_7329; // @[Mux.scala 31:69:@3957.4]
  assign _T_7331 = _T_7330[0]; // @[OneHot.scala 66:30:@3958.4]
  assign _T_7332 = _T_7330[1]; // @[OneHot.scala 66:30:@3959.4]
  assign _T_7333 = _T_7330[2]; // @[OneHot.scala 66:30:@3960.4]
  assign _T_7334 = _T_7330[3]; // @[OneHot.scala 66:30:@3961.4]
  assign _T_7335 = _T_7330[4]; // @[OneHot.scala 66:30:@3962.4]
  assign _T_7336 = _T_7330[5]; // @[OneHot.scala 66:30:@3963.4]
  assign _T_7337 = _T_7330[6]; // @[OneHot.scala 66:30:@3964.4]
  assign _T_7338 = _T_7330[7]; // @[OneHot.scala 66:30:@3965.4]
  assign _T_7339 = _T_7330[8]; // @[OneHot.scala 66:30:@3966.4]
  assign _T_7340 = _T_7330[9]; // @[OneHot.scala 66:30:@3967.4]
  assign _T_7341 = _T_7330[10]; // @[OneHot.scala 66:30:@3968.4]
  assign _T_7342 = _T_7330[11]; // @[OneHot.scala 66:30:@3969.4]
  assign _T_7343 = _T_7330[12]; // @[OneHot.scala 66:30:@3970.4]
  assign _T_7344 = _T_7330[13]; // @[OneHot.scala 66:30:@3971.4]
  assign _T_7345 = _T_7330[14]; // @[OneHot.scala 66:30:@3972.4]
  assign _T_7346 = _T_7330[15]; // @[OneHot.scala 66:30:@3973.4]
  assign _T_7411 = {_T_6258,_T_6257,_T_6256,_T_6255,_T_6254,_T_6253,_T_6252,_T_6251}; // @[Mux.scala 19:72:@3997.4]
  assign _T_7419 = {_T_6266,_T_6265,_T_6264,_T_6263,_T_6262,_T_6261,_T_6260,_T_6259,_T_7411}; // @[Mux.scala 19:72:@4005.4]
  assign _T_7421 = _T_4521 ? _T_7419 : 16'h0; // @[Mux.scala 19:72:@4006.4]
  assign _T_7428 = {_T_6329,_T_6328,_T_6327,_T_6326,_T_6325,_T_6324,_T_6323,_T_6338}; // @[Mux.scala 19:72:@4013.4]
  assign _T_7436 = {_T_6337,_T_6336,_T_6335,_T_6334,_T_6333,_T_6332,_T_6331,_T_6330,_T_7428}; // @[Mux.scala 19:72:@4021.4]
  assign _T_7438 = _T_4522 ? _T_7436 : 16'h0; // @[Mux.scala 19:72:@4022.4]
  assign _T_7445 = {_T_6400,_T_6399,_T_6398,_T_6397,_T_6396,_T_6395,_T_6410,_T_6409}; // @[Mux.scala 19:72:@4029.4]
  assign _T_7453 = {_T_6408,_T_6407,_T_6406,_T_6405,_T_6404,_T_6403,_T_6402,_T_6401,_T_7445}; // @[Mux.scala 19:72:@4037.4]
  assign _T_7455 = _T_4523 ? _T_7453 : 16'h0; // @[Mux.scala 19:72:@4038.4]
  assign _T_7462 = {_T_6471,_T_6470,_T_6469,_T_6468,_T_6467,_T_6482,_T_6481,_T_6480}; // @[Mux.scala 19:72:@4045.4]
  assign _T_7470 = {_T_6479,_T_6478,_T_6477,_T_6476,_T_6475,_T_6474,_T_6473,_T_6472,_T_7462}; // @[Mux.scala 19:72:@4053.4]
  assign _T_7472 = _T_4524 ? _T_7470 : 16'h0; // @[Mux.scala 19:72:@4054.4]
  assign _T_7479 = {_T_6542,_T_6541,_T_6540,_T_6539,_T_6554,_T_6553,_T_6552,_T_6551}; // @[Mux.scala 19:72:@4061.4]
  assign _T_7487 = {_T_6550,_T_6549,_T_6548,_T_6547,_T_6546,_T_6545,_T_6544,_T_6543,_T_7479}; // @[Mux.scala 19:72:@4069.4]
  assign _T_7489 = _T_4525 ? _T_7487 : 16'h0; // @[Mux.scala 19:72:@4070.4]
  assign _T_7496 = {_T_6613,_T_6612,_T_6611,_T_6626,_T_6625,_T_6624,_T_6623,_T_6622}; // @[Mux.scala 19:72:@4077.4]
  assign _T_7504 = {_T_6621,_T_6620,_T_6619,_T_6618,_T_6617,_T_6616,_T_6615,_T_6614,_T_7496}; // @[Mux.scala 19:72:@4085.4]
  assign _T_7506 = _T_4526 ? _T_7504 : 16'h0; // @[Mux.scala 19:72:@4086.4]
  assign _T_7513 = {_T_6684,_T_6683,_T_6698,_T_6697,_T_6696,_T_6695,_T_6694,_T_6693}; // @[Mux.scala 19:72:@4093.4]
  assign _T_7521 = {_T_6692,_T_6691,_T_6690,_T_6689,_T_6688,_T_6687,_T_6686,_T_6685,_T_7513}; // @[Mux.scala 19:72:@4101.4]
  assign _T_7523 = _T_4527 ? _T_7521 : 16'h0; // @[Mux.scala 19:72:@4102.4]
  assign _T_7530 = {_T_6755,_T_6770,_T_6769,_T_6768,_T_6767,_T_6766,_T_6765,_T_6764}; // @[Mux.scala 19:72:@4109.4]
  assign _T_7538 = {_T_6763,_T_6762,_T_6761,_T_6760,_T_6759,_T_6758,_T_6757,_T_6756,_T_7530}; // @[Mux.scala 19:72:@4117.4]
  assign _T_7540 = _T_4528 ? _T_7538 : 16'h0; // @[Mux.scala 19:72:@4118.4]
  assign _T_7547 = {_T_6842,_T_6841,_T_6840,_T_6839,_T_6838,_T_6837,_T_6836,_T_6835}; // @[Mux.scala 19:72:@4125.4]
  assign _T_7555 = {_T_6834,_T_6833,_T_6832,_T_6831,_T_6830,_T_6829,_T_6828,_T_6827,_T_7547}; // @[Mux.scala 19:72:@4133.4]
  assign _T_7557 = _T_4529 ? _T_7555 : 16'h0; // @[Mux.scala 19:72:@4134.4]
  assign _T_7564 = {_T_6913,_T_6912,_T_6911,_T_6910,_T_6909,_T_6908,_T_6907,_T_6906}; // @[Mux.scala 19:72:@4141.4]
  assign _T_7572 = {_T_6905,_T_6904,_T_6903,_T_6902,_T_6901,_T_6900,_T_6899,_T_6914,_T_7564}; // @[Mux.scala 19:72:@4149.4]
  assign _T_7574 = _T_4530 ? _T_7572 : 16'h0; // @[Mux.scala 19:72:@4150.4]
  assign _T_7581 = {_T_6984,_T_6983,_T_6982,_T_6981,_T_6980,_T_6979,_T_6978,_T_6977}; // @[Mux.scala 19:72:@4157.4]
  assign _T_7589 = {_T_6976,_T_6975,_T_6974,_T_6973,_T_6972,_T_6971,_T_6986,_T_6985,_T_7581}; // @[Mux.scala 19:72:@4165.4]
  assign _T_7591 = _T_4531 ? _T_7589 : 16'h0; // @[Mux.scala 19:72:@4166.4]
  assign _T_7598 = {_T_7055,_T_7054,_T_7053,_T_7052,_T_7051,_T_7050,_T_7049,_T_7048}; // @[Mux.scala 19:72:@4173.4]
  assign _T_7606 = {_T_7047,_T_7046,_T_7045,_T_7044,_T_7043,_T_7058,_T_7057,_T_7056,_T_7598}; // @[Mux.scala 19:72:@4181.4]
  assign _T_7608 = _T_4532 ? _T_7606 : 16'h0; // @[Mux.scala 19:72:@4182.4]
  assign _T_7615 = {_T_7126,_T_7125,_T_7124,_T_7123,_T_7122,_T_7121,_T_7120,_T_7119}; // @[Mux.scala 19:72:@4189.4]
  assign _T_7623 = {_T_7118,_T_7117,_T_7116,_T_7115,_T_7130,_T_7129,_T_7128,_T_7127,_T_7615}; // @[Mux.scala 19:72:@4197.4]
  assign _T_7625 = _T_4533 ? _T_7623 : 16'h0; // @[Mux.scala 19:72:@4198.4]
  assign _T_7632 = {_T_7197,_T_7196,_T_7195,_T_7194,_T_7193,_T_7192,_T_7191,_T_7190}; // @[Mux.scala 19:72:@4205.4]
  assign _T_7640 = {_T_7189,_T_7188,_T_7187,_T_7202,_T_7201,_T_7200,_T_7199,_T_7198,_T_7632}; // @[Mux.scala 19:72:@4213.4]
  assign _T_7642 = _T_4534 ? _T_7640 : 16'h0; // @[Mux.scala 19:72:@4214.4]
  assign _T_7649 = {_T_7268,_T_7267,_T_7266,_T_7265,_T_7264,_T_7263,_T_7262,_T_7261}; // @[Mux.scala 19:72:@4221.4]
  assign _T_7657 = {_T_7260,_T_7259,_T_7274,_T_7273,_T_7272,_T_7271,_T_7270,_T_7269,_T_7649}; // @[Mux.scala 19:72:@4229.4]
  assign _T_7659 = _T_4535 ? _T_7657 : 16'h0; // @[Mux.scala 19:72:@4230.4]
  assign _T_7666 = {_T_7339,_T_7338,_T_7337,_T_7336,_T_7335,_T_7334,_T_7333,_T_7332}; // @[Mux.scala 19:72:@4237.4]
  assign _T_7674 = {_T_7331,_T_7346,_T_7345,_T_7344,_T_7343,_T_7342,_T_7341,_T_7340,_T_7666}; // @[Mux.scala 19:72:@4245.4]
  assign _T_7676 = _T_4536 ? _T_7674 : 16'h0; // @[Mux.scala 19:72:@4246.4]
  assign _T_7677 = _T_7421 | _T_7438; // @[Mux.scala 19:72:@4247.4]
  assign _T_7678 = _T_7677 | _T_7455; // @[Mux.scala 19:72:@4248.4]
  assign _T_7679 = _T_7678 | _T_7472; // @[Mux.scala 19:72:@4249.4]
  assign _T_7680 = _T_7679 | _T_7489; // @[Mux.scala 19:72:@4250.4]
  assign _T_7681 = _T_7680 | _T_7506; // @[Mux.scala 19:72:@4251.4]
  assign _T_7682 = _T_7681 | _T_7523; // @[Mux.scala 19:72:@4252.4]
  assign _T_7683 = _T_7682 | _T_7540; // @[Mux.scala 19:72:@4253.4]
  assign _T_7684 = _T_7683 | _T_7557; // @[Mux.scala 19:72:@4254.4]
  assign _T_7685 = _T_7684 | _T_7574; // @[Mux.scala 19:72:@4255.4]
  assign _T_7686 = _T_7685 | _T_7591; // @[Mux.scala 19:72:@4256.4]
  assign _T_7687 = _T_7686 | _T_7608; // @[Mux.scala 19:72:@4257.4]
  assign _T_7688 = _T_7687 | _T_7625; // @[Mux.scala 19:72:@4258.4]
  assign _T_7689 = _T_7688 | _T_7642; // @[Mux.scala 19:72:@4259.4]
  assign _T_7690 = _T_7689 | _T_7659; // @[Mux.scala 19:72:@4260.4]
  assign _T_7691 = _T_7690 | _T_7676; // @[Mux.scala 19:72:@4261.4]
  assign inputDataPriorityPorts_0_0 = _T_7691[0]; // @[Mux.scala 19:72:@4265.4]
  assign inputDataPriorityPorts_0_1 = _T_7691[1]; // @[Mux.scala 19:72:@4267.4]
  assign inputDataPriorityPorts_0_2 = _T_7691[2]; // @[Mux.scala 19:72:@4269.4]
  assign inputDataPriorityPorts_0_3 = _T_7691[3]; // @[Mux.scala 19:72:@4271.4]
  assign inputDataPriorityPorts_0_4 = _T_7691[4]; // @[Mux.scala 19:72:@4273.4]
  assign inputDataPriorityPorts_0_5 = _T_7691[5]; // @[Mux.scala 19:72:@4275.4]
  assign inputDataPriorityPorts_0_6 = _T_7691[6]; // @[Mux.scala 19:72:@4277.4]
  assign inputDataPriorityPorts_0_7 = _T_7691[7]; // @[Mux.scala 19:72:@4279.4]
  assign inputDataPriorityPorts_0_8 = _T_7691[8]; // @[Mux.scala 19:72:@4281.4]
  assign inputDataPriorityPorts_0_9 = _T_7691[9]; // @[Mux.scala 19:72:@4283.4]
  assign inputDataPriorityPorts_0_10 = _T_7691[10]; // @[Mux.scala 19:72:@4285.4]
  assign inputDataPriorityPorts_0_11 = _T_7691[11]; // @[Mux.scala 19:72:@4287.4]
  assign inputDataPriorityPorts_0_12 = _T_7691[12]; // @[Mux.scala 19:72:@4289.4]
  assign inputDataPriorityPorts_0_13 = _T_7691[13]; // @[Mux.scala 19:72:@4291.4]
  assign inputDataPriorityPorts_0_14 = _T_7691[14]; // @[Mux.scala 19:72:@4293.4]
  assign inputDataPriorityPorts_0_15 = _T_7691[15]; // @[Mux.scala 19:72:@4295.4]
  assign _T_7835 = portQ_0 & _T_4378; // @[StoreQueue.scala 192:88:@4314.4]
  assign _T_7838 = portQ_1 & _T_4381; // @[StoreQueue.scala 192:88:@4316.4]
  assign _T_7841 = portQ_2 & _T_4384; // @[StoreQueue.scala 192:88:@4318.4]
  assign _T_7844 = portQ_3 & _T_4387; // @[StoreQueue.scala 192:88:@4320.4]
  assign _T_7847 = portQ_4 & _T_4390; // @[StoreQueue.scala 192:88:@4322.4]
  assign _T_7850 = portQ_5 & _T_4393; // @[StoreQueue.scala 192:88:@4324.4]
  assign _T_7853 = portQ_6 & _T_4396; // @[StoreQueue.scala 192:88:@4326.4]
  assign _T_7856 = portQ_7 & _T_4399; // @[StoreQueue.scala 192:88:@4328.4]
  assign _T_7859 = portQ_8 & _T_4402; // @[StoreQueue.scala 192:88:@4330.4]
  assign _T_7862 = portQ_9 & _T_4405; // @[StoreQueue.scala 192:88:@4332.4]
  assign _T_7865 = portQ_10 & _T_4408; // @[StoreQueue.scala 192:88:@4334.4]
  assign _T_7868 = portQ_11 & _T_4411; // @[StoreQueue.scala 192:88:@4336.4]
  assign _T_7871 = portQ_12 & _T_4414; // @[StoreQueue.scala 192:88:@4338.4]
  assign _T_7874 = portQ_13 & _T_4417; // @[StoreQueue.scala 192:88:@4340.4]
  assign _T_7877 = portQ_14 & _T_4420; // @[StoreQueue.scala 192:88:@4342.4]
  assign _T_7880 = portQ_15 & _T_4423; // @[StoreQueue.scala 192:88:@4344.4]
  assign _T_7905 = portQ_0 & _T_4448; // @[StoreQueue.scala 193:88:@4363.4]
  assign _T_7908 = portQ_1 & _T_4451; // @[StoreQueue.scala 193:88:@4365.4]
  assign _T_7911 = portQ_2 & _T_4454; // @[StoreQueue.scala 193:88:@4367.4]
  assign _T_7914 = portQ_3 & _T_4457; // @[StoreQueue.scala 193:88:@4369.4]
  assign _T_7917 = portQ_4 & _T_4460; // @[StoreQueue.scala 193:88:@4371.4]
  assign _T_7920 = portQ_5 & _T_4463; // @[StoreQueue.scala 193:88:@4373.4]
  assign _T_7923 = portQ_6 & _T_4466; // @[StoreQueue.scala 193:88:@4375.4]
  assign _T_7926 = portQ_7 & _T_4469; // @[StoreQueue.scala 193:88:@4377.4]
  assign _T_7929 = portQ_8 & _T_4472; // @[StoreQueue.scala 193:88:@4379.4]
  assign _T_7932 = portQ_9 & _T_4475; // @[StoreQueue.scala 193:88:@4381.4]
  assign _T_7935 = portQ_10 & _T_4478; // @[StoreQueue.scala 193:88:@4383.4]
  assign _T_7938 = portQ_11 & _T_4481; // @[StoreQueue.scala 193:88:@4385.4]
  assign _T_7941 = portQ_12 & _T_4484; // @[StoreQueue.scala 193:88:@4387.4]
  assign _T_7944 = portQ_13 & _T_4487; // @[StoreQueue.scala 193:88:@4389.4]
  assign _T_7947 = portQ_14 & _T_4490; // @[StoreQueue.scala 193:88:@4391.4]
  assign _T_7950 = portQ_15 & _T_4493; // @[StoreQueue.scala 193:88:@4393.4]
  assign _T_8033 = _T_7880 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4447.4]
  assign _T_8034 = _T_7877 ? 16'h4000 : _T_8033; // @[Mux.scala 31:69:@4448.4]
  assign _T_8035 = _T_7874 ? 16'h2000 : _T_8034; // @[Mux.scala 31:69:@4449.4]
  assign _T_8036 = _T_7871 ? 16'h1000 : _T_8035; // @[Mux.scala 31:69:@4450.4]
  assign _T_8037 = _T_7868 ? 16'h800 : _T_8036; // @[Mux.scala 31:69:@4451.4]
  assign _T_8038 = _T_7865 ? 16'h400 : _T_8037; // @[Mux.scala 31:69:@4452.4]
  assign _T_8039 = _T_7862 ? 16'h200 : _T_8038; // @[Mux.scala 31:69:@4453.4]
  assign _T_8040 = _T_7859 ? 16'h100 : _T_8039; // @[Mux.scala 31:69:@4454.4]
  assign _T_8041 = _T_7856 ? 16'h80 : _T_8040; // @[Mux.scala 31:69:@4455.4]
  assign _T_8042 = _T_7853 ? 16'h40 : _T_8041; // @[Mux.scala 31:69:@4456.4]
  assign _T_8043 = _T_7850 ? 16'h20 : _T_8042; // @[Mux.scala 31:69:@4457.4]
  assign _T_8044 = _T_7847 ? 16'h10 : _T_8043; // @[Mux.scala 31:69:@4458.4]
  assign _T_8045 = _T_7844 ? 16'h8 : _T_8044; // @[Mux.scala 31:69:@4459.4]
  assign _T_8046 = _T_7841 ? 16'h4 : _T_8045; // @[Mux.scala 31:69:@4460.4]
  assign _T_8047 = _T_7838 ? 16'h2 : _T_8046; // @[Mux.scala 31:69:@4461.4]
  assign _T_8048 = _T_7835 ? 16'h1 : _T_8047; // @[Mux.scala 31:69:@4462.4]
  assign _T_8049 = _T_8048[0]; // @[OneHot.scala 66:30:@4463.4]
  assign _T_8050 = _T_8048[1]; // @[OneHot.scala 66:30:@4464.4]
  assign _T_8051 = _T_8048[2]; // @[OneHot.scala 66:30:@4465.4]
  assign _T_8052 = _T_8048[3]; // @[OneHot.scala 66:30:@4466.4]
  assign _T_8053 = _T_8048[4]; // @[OneHot.scala 66:30:@4467.4]
  assign _T_8054 = _T_8048[5]; // @[OneHot.scala 66:30:@4468.4]
  assign _T_8055 = _T_8048[6]; // @[OneHot.scala 66:30:@4469.4]
  assign _T_8056 = _T_8048[7]; // @[OneHot.scala 66:30:@4470.4]
  assign _T_8057 = _T_8048[8]; // @[OneHot.scala 66:30:@4471.4]
  assign _T_8058 = _T_8048[9]; // @[OneHot.scala 66:30:@4472.4]
  assign _T_8059 = _T_8048[10]; // @[OneHot.scala 66:30:@4473.4]
  assign _T_8060 = _T_8048[11]; // @[OneHot.scala 66:30:@4474.4]
  assign _T_8061 = _T_8048[12]; // @[OneHot.scala 66:30:@4475.4]
  assign _T_8062 = _T_8048[13]; // @[OneHot.scala 66:30:@4476.4]
  assign _T_8063 = _T_8048[14]; // @[OneHot.scala 66:30:@4477.4]
  assign _T_8064 = _T_8048[15]; // @[OneHot.scala 66:30:@4478.4]
  assign _T_8105 = _T_7835 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4496.4]
  assign _T_8106 = _T_7880 ? 16'h4000 : _T_8105; // @[Mux.scala 31:69:@4497.4]
  assign _T_8107 = _T_7877 ? 16'h2000 : _T_8106; // @[Mux.scala 31:69:@4498.4]
  assign _T_8108 = _T_7874 ? 16'h1000 : _T_8107; // @[Mux.scala 31:69:@4499.4]
  assign _T_8109 = _T_7871 ? 16'h800 : _T_8108; // @[Mux.scala 31:69:@4500.4]
  assign _T_8110 = _T_7868 ? 16'h400 : _T_8109; // @[Mux.scala 31:69:@4501.4]
  assign _T_8111 = _T_7865 ? 16'h200 : _T_8110; // @[Mux.scala 31:69:@4502.4]
  assign _T_8112 = _T_7862 ? 16'h100 : _T_8111; // @[Mux.scala 31:69:@4503.4]
  assign _T_8113 = _T_7859 ? 16'h80 : _T_8112; // @[Mux.scala 31:69:@4504.4]
  assign _T_8114 = _T_7856 ? 16'h40 : _T_8113; // @[Mux.scala 31:69:@4505.4]
  assign _T_8115 = _T_7853 ? 16'h20 : _T_8114; // @[Mux.scala 31:69:@4506.4]
  assign _T_8116 = _T_7850 ? 16'h10 : _T_8115; // @[Mux.scala 31:69:@4507.4]
  assign _T_8117 = _T_7847 ? 16'h8 : _T_8116; // @[Mux.scala 31:69:@4508.4]
  assign _T_8118 = _T_7844 ? 16'h4 : _T_8117; // @[Mux.scala 31:69:@4509.4]
  assign _T_8119 = _T_7841 ? 16'h2 : _T_8118; // @[Mux.scala 31:69:@4510.4]
  assign _T_8120 = _T_7838 ? 16'h1 : _T_8119; // @[Mux.scala 31:69:@4511.4]
  assign _T_8121 = _T_8120[0]; // @[OneHot.scala 66:30:@4512.4]
  assign _T_8122 = _T_8120[1]; // @[OneHot.scala 66:30:@4513.4]
  assign _T_8123 = _T_8120[2]; // @[OneHot.scala 66:30:@4514.4]
  assign _T_8124 = _T_8120[3]; // @[OneHot.scala 66:30:@4515.4]
  assign _T_8125 = _T_8120[4]; // @[OneHot.scala 66:30:@4516.4]
  assign _T_8126 = _T_8120[5]; // @[OneHot.scala 66:30:@4517.4]
  assign _T_8127 = _T_8120[6]; // @[OneHot.scala 66:30:@4518.4]
  assign _T_8128 = _T_8120[7]; // @[OneHot.scala 66:30:@4519.4]
  assign _T_8129 = _T_8120[8]; // @[OneHot.scala 66:30:@4520.4]
  assign _T_8130 = _T_8120[9]; // @[OneHot.scala 66:30:@4521.4]
  assign _T_8131 = _T_8120[10]; // @[OneHot.scala 66:30:@4522.4]
  assign _T_8132 = _T_8120[11]; // @[OneHot.scala 66:30:@4523.4]
  assign _T_8133 = _T_8120[12]; // @[OneHot.scala 66:30:@4524.4]
  assign _T_8134 = _T_8120[13]; // @[OneHot.scala 66:30:@4525.4]
  assign _T_8135 = _T_8120[14]; // @[OneHot.scala 66:30:@4526.4]
  assign _T_8136 = _T_8120[15]; // @[OneHot.scala 66:30:@4527.4]
  assign _T_8177 = _T_7838 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4545.4]
  assign _T_8178 = _T_7835 ? 16'h4000 : _T_8177; // @[Mux.scala 31:69:@4546.4]
  assign _T_8179 = _T_7880 ? 16'h2000 : _T_8178; // @[Mux.scala 31:69:@4547.4]
  assign _T_8180 = _T_7877 ? 16'h1000 : _T_8179; // @[Mux.scala 31:69:@4548.4]
  assign _T_8181 = _T_7874 ? 16'h800 : _T_8180; // @[Mux.scala 31:69:@4549.4]
  assign _T_8182 = _T_7871 ? 16'h400 : _T_8181; // @[Mux.scala 31:69:@4550.4]
  assign _T_8183 = _T_7868 ? 16'h200 : _T_8182; // @[Mux.scala 31:69:@4551.4]
  assign _T_8184 = _T_7865 ? 16'h100 : _T_8183; // @[Mux.scala 31:69:@4552.4]
  assign _T_8185 = _T_7862 ? 16'h80 : _T_8184; // @[Mux.scala 31:69:@4553.4]
  assign _T_8186 = _T_7859 ? 16'h40 : _T_8185; // @[Mux.scala 31:69:@4554.4]
  assign _T_8187 = _T_7856 ? 16'h20 : _T_8186; // @[Mux.scala 31:69:@4555.4]
  assign _T_8188 = _T_7853 ? 16'h10 : _T_8187; // @[Mux.scala 31:69:@4556.4]
  assign _T_8189 = _T_7850 ? 16'h8 : _T_8188; // @[Mux.scala 31:69:@4557.4]
  assign _T_8190 = _T_7847 ? 16'h4 : _T_8189; // @[Mux.scala 31:69:@4558.4]
  assign _T_8191 = _T_7844 ? 16'h2 : _T_8190; // @[Mux.scala 31:69:@4559.4]
  assign _T_8192 = _T_7841 ? 16'h1 : _T_8191; // @[Mux.scala 31:69:@4560.4]
  assign _T_8193 = _T_8192[0]; // @[OneHot.scala 66:30:@4561.4]
  assign _T_8194 = _T_8192[1]; // @[OneHot.scala 66:30:@4562.4]
  assign _T_8195 = _T_8192[2]; // @[OneHot.scala 66:30:@4563.4]
  assign _T_8196 = _T_8192[3]; // @[OneHot.scala 66:30:@4564.4]
  assign _T_8197 = _T_8192[4]; // @[OneHot.scala 66:30:@4565.4]
  assign _T_8198 = _T_8192[5]; // @[OneHot.scala 66:30:@4566.4]
  assign _T_8199 = _T_8192[6]; // @[OneHot.scala 66:30:@4567.4]
  assign _T_8200 = _T_8192[7]; // @[OneHot.scala 66:30:@4568.4]
  assign _T_8201 = _T_8192[8]; // @[OneHot.scala 66:30:@4569.4]
  assign _T_8202 = _T_8192[9]; // @[OneHot.scala 66:30:@4570.4]
  assign _T_8203 = _T_8192[10]; // @[OneHot.scala 66:30:@4571.4]
  assign _T_8204 = _T_8192[11]; // @[OneHot.scala 66:30:@4572.4]
  assign _T_8205 = _T_8192[12]; // @[OneHot.scala 66:30:@4573.4]
  assign _T_8206 = _T_8192[13]; // @[OneHot.scala 66:30:@4574.4]
  assign _T_8207 = _T_8192[14]; // @[OneHot.scala 66:30:@4575.4]
  assign _T_8208 = _T_8192[15]; // @[OneHot.scala 66:30:@4576.4]
  assign _T_8249 = _T_7841 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4594.4]
  assign _T_8250 = _T_7838 ? 16'h4000 : _T_8249; // @[Mux.scala 31:69:@4595.4]
  assign _T_8251 = _T_7835 ? 16'h2000 : _T_8250; // @[Mux.scala 31:69:@4596.4]
  assign _T_8252 = _T_7880 ? 16'h1000 : _T_8251; // @[Mux.scala 31:69:@4597.4]
  assign _T_8253 = _T_7877 ? 16'h800 : _T_8252; // @[Mux.scala 31:69:@4598.4]
  assign _T_8254 = _T_7874 ? 16'h400 : _T_8253; // @[Mux.scala 31:69:@4599.4]
  assign _T_8255 = _T_7871 ? 16'h200 : _T_8254; // @[Mux.scala 31:69:@4600.4]
  assign _T_8256 = _T_7868 ? 16'h100 : _T_8255; // @[Mux.scala 31:69:@4601.4]
  assign _T_8257 = _T_7865 ? 16'h80 : _T_8256; // @[Mux.scala 31:69:@4602.4]
  assign _T_8258 = _T_7862 ? 16'h40 : _T_8257; // @[Mux.scala 31:69:@4603.4]
  assign _T_8259 = _T_7859 ? 16'h20 : _T_8258; // @[Mux.scala 31:69:@4604.4]
  assign _T_8260 = _T_7856 ? 16'h10 : _T_8259; // @[Mux.scala 31:69:@4605.4]
  assign _T_8261 = _T_7853 ? 16'h8 : _T_8260; // @[Mux.scala 31:69:@4606.4]
  assign _T_8262 = _T_7850 ? 16'h4 : _T_8261; // @[Mux.scala 31:69:@4607.4]
  assign _T_8263 = _T_7847 ? 16'h2 : _T_8262; // @[Mux.scala 31:69:@4608.4]
  assign _T_8264 = _T_7844 ? 16'h1 : _T_8263; // @[Mux.scala 31:69:@4609.4]
  assign _T_8265 = _T_8264[0]; // @[OneHot.scala 66:30:@4610.4]
  assign _T_8266 = _T_8264[1]; // @[OneHot.scala 66:30:@4611.4]
  assign _T_8267 = _T_8264[2]; // @[OneHot.scala 66:30:@4612.4]
  assign _T_8268 = _T_8264[3]; // @[OneHot.scala 66:30:@4613.4]
  assign _T_8269 = _T_8264[4]; // @[OneHot.scala 66:30:@4614.4]
  assign _T_8270 = _T_8264[5]; // @[OneHot.scala 66:30:@4615.4]
  assign _T_8271 = _T_8264[6]; // @[OneHot.scala 66:30:@4616.4]
  assign _T_8272 = _T_8264[7]; // @[OneHot.scala 66:30:@4617.4]
  assign _T_8273 = _T_8264[8]; // @[OneHot.scala 66:30:@4618.4]
  assign _T_8274 = _T_8264[9]; // @[OneHot.scala 66:30:@4619.4]
  assign _T_8275 = _T_8264[10]; // @[OneHot.scala 66:30:@4620.4]
  assign _T_8276 = _T_8264[11]; // @[OneHot.scala 66:30:@4621.4]
  assign _T_8277 = _T_8264[12]; // @[OneHot.scala 66:30:@4622.4]
  assign _T_8278 = _T_8264[13]; // @[OneHot.scala 66:30:@4623.4]
  assign _T_8279 = _T_8264[14]; // @[OneHot.scala 66:30:@4624.4]
  assign _T_8280 = _T_8264[15]; // @[OneHot.scala 66:30:@4625.4]
  assign _T_8321 = _T_7844 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4643.4]
  assign _T_8322 = _T_7841 ? 16'h4000 : _T_8321; // @[Mux.scala 31:69:@4644.4]
  assign _T_8323 = _T_7838 ? 16'h2000 : _T_8322; // @[Mux.scala 31:69:@4645.4]
  assign _T_8324 = _T_7835 ? 16'h1000 : _T_8323; // @[Mux.scala 31:69:@4646.4]
  assign _T_8325 = _T_7880 ? 16'h800 : _T_8324; // @[Mux.scala 31:69:@4647.4]
  assign _T_8326 = _T_7877 ? 16'h400 : _T_8325; // @[Mux.scala 31:69:@4648.4]
  assign _T_8327 = _T_7874 ? 16'h200 : _T_8326; // @[Mux.scala 31:69:@4649.4]
  assign _T_8328 = _T_7871 ? 16'h100 : _T_8327; // @[Mux.scala 31:69:@4650.4]
  assign _T_8329 = _T_7868 ? 16'h80 : _T_8328; // @[Mux.scala 31:69:@4651.4]
  assign _T_8330 = _T_7865 ? 16'h40 : _T_8329; // @[Mux.scala 31:69:@4652.4]
  assign _T_8331 = _T_7862 ? 16'h20 : _T_8330; // @[Mux.scala 31:69:@4653.4]
  assign _T_8332 = _T_7859 ? 16'h10 : _T_8331; // @[Mux.scala 31:69:@4654.4]
  assign _T_8333 = _T_7856 ? 16'h8 : _T_8332; // @[Mux.scala 31:69:@4655.4]
  assign _T_8334 = _T_7853 ? 16'h4 : _T_8333; // @[Mux.scala 31:69:@4656.4]
  assign _T_8335 = _T_7850 ? 16'h2 : _T_8334; // @[Mux.scala 31:69:@4657.4]
  assign _T_8336 = _T_7847 ? 16'h1 : _T_8335; // @[Mux.scala 31:69:@4658.4]
  assign _T_8337 = _T_8336[0]; // @[OneHot.scala 66:30:@4659.4]
  assign _T_8338 = _T_8336[1]; // @[OneHot.scala 66:30:@4660.4]
  assign _T_8339 = _T_8336[2]; // @[OneHot.scala 66:30:@4661.4]
  assign _T_8340 = _T_8336[3]; // @[OneHot.scala 66:30:@4662.4]
  assign _T_8341 = _T_8336[4]; // @[OneHot.scala 66:30:@4663.4]
  assign _T_8342 = _T_8336[5]; // @[OneHot.scala 66:30:@4664.4]
  assign _T_8343 = _T_8336[6]; // @[OneHot.scala 66:30:@4665.4]
  assign _T_8344 = _T_8336[7]; // @[OneHot.scala 66:30:@4666.4]
  assign _T_8345 = _T_8336[8]; // @[OneHot.scala 66:30:@4667.4]
  assign _T_8346 = _T_8336[9]; // @[OneHot.scala 66:30:@4668.4]
  assign _T_8347 = _T_8336[10]; // @[OneHot.scala 66:30:@4669.4]
  assign _T_8348 = _T_8336[11]; // @[OneHot.scala 66:30:@4670.4]
  assign _T_8349 = _T_8336[12]; // @[OneHot.scala 66:30:@4671.4]
  assign _T_8350 = _T_8336[13]; // @[OneHot.scala 66:30:@4672.4]
  assign _T_8351 = _T_8336[14]; // @[OneHot.scala 66:30:@4673.4]
  assign _T_8352 = _T_8336[15]; // @[OneHot.scala 66:30:@4674.4]
  assign _T_8393 = _T_7847 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4692.4]
  assign _T_8394 = _T_7844 ? 16'h4000 : _T_8393; // @[Mux.scala 31:69:@4693.4]
  assign _T_8395 = _T_7841 ? 16'h2000 : _T_8394; // @[Mux.scala 31:69:@4694.4]
  assign _T_8396 = _T_7838 ? 16'h1000 : _T_8395; // @[Mux.scala 31:69:@4695.4]
  assign _T_8397 = _T_7835 ? 16'h800 : _T_8396; // @[Mux.scala 31:69:@4696.4]
  assign _T_8398 = _T_7880 ? 16'h400 : _T_8397; // @[Mux.scala 31:69:@4697.4]
  assign _T_8399 = _T_7877 ? 16'h200 : _T_8398; // @[Mux.scala 31:69:@4698.4]
  assign _T_8400 = _T_7874 ? 16'h100 : _T_8399; // @[Mux.scala 31:69:@4699.4]
  assign _T_8401 = _T_7871 ? 16'h80 : _T_8400; // @[Mux.scala 31:69:@4700.4]
  assign _T_8402 = _T_7868 ? 16'h40 : _T_8401; // @[Mux.scala 31:69:@4701.4]
  assign _T_8403 = _T_7865 ? 16'h20 : _T_8402; // @[Mux.scala 31:69:@4702.4]
  assign _T_8404 = _T_7862 ? 16'h10 : _T_8403; // @[Mux.scala 31:69:@4703.4]
  assign _T_8405 = _T_7859 ? 16'h8 : _T_8404; // @[Mux.scala 31:69:@4704.4]
  assign _T_8406 = _T_7856 ? 16'h4 : _T_8405; // @[Mux.scala 31:69:@4705.4]
  assign _T_8407 = _T_7853 ? 16'h2 : _T_8406; // @[Mux.scala 31:69:@4706.4]
  assign _T_8408 = _T_7850 ? 16'h1 : _T_8407; // @[Mux.scala 31:69:@4707.4]
  assign _T_8409 = _T_8408[0]; // @[OneHot.scala 66:30:@4708.4]
  assign _T_8410 = _T_8408[1]; // @[OneHot.scala 66:30:@4709.4]
  assign _T_8411 = _T_8408[2]; // @[OneHot.scala 66:30:@4710.4]
  assign _T_8412 = _T_8408[3]; // @[OneHot.scala 66:30:@4711.4]
  assign _T_8413 = _T_8408[4]; // @[OneHot.scala 66:30:@4712.4]
  assign _T_8414 = _T_8408[5]; // @[OneHot.scala 66:30:@4713.4]
  assign _T_8415 = _T_8408[6]; // @[OneHot.scala 66:30:@4714.4]
  assign _T_8416 = _T_8408[7]; // @[OneHot.scala 66:30:@4715.4]
  assign _T_8417 = _T_8408[8]; // @[OneHot.scala 66:30:@4716.4]
  assign _T_8418 = _T_8408[9]; // @[OneHot.scala 66:30:@4717.4]
  assign _T_8419 = _T_8408[10]; // @[OneHot.scala 66:30:@4718.4]
  assign _T_8420 = _T_8408[11]; // @[OneHot.scala 66:30:@4719.4]
  assign _T_8421 = _T_8408[12]; // @[OneHot.scala 66:30:@4720.4]
  assign _T_8422 = _T_8408[13]; // @[OneHot.scala 66:30:@4721.4]
  assign _T_8423 = _T_8408[14]; // @[OneHot.scala 66:30:@4722.4]
  assign _T_8424 = _T_8408[15]; // @[OneHot.scala 66:30:@4723.4]
  assign _T_8465 = _T_7850 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4741.4]
  assign _T_8466 = _T_7847 ? 16'h4000 : _T_8465; // @[Mux.scala 31:69:@4742.4]
  assign _T_8467 = _T_7844 ? 16'h2000 : _T_8466; // @[Mux.scala 31:69:@4743.4]
  assign _T_8468 = _T_7841 ? 16'h1000 : _T_8467; // @[Mux.scala 31:69:@4744.4]
  assign _T_8469 = _T_7838 ? 16'h800 : _T_8468; // @[Mux.scala 31:69:@4745.4]
  assign _T_8470 = _T_7835 ? 16'h400 : _T_8469; // @[Mux.scala 31:69:@4746.4]
  assign _T_8471 = _T_7880 ? 16'h200 : _T_8470; // @[Mux.scala 31:69:@4747.4]
  assign _T_8472 = _T_7877 ? 16'h100 : _T_8471; // @[Mux.scala 31:69:@4748.4]
  assign _T_8473 = _T_7874 ? 16'h80 : _T_8472; // @[Mux.scala 31:69:@4749.4]
  assign _T_8474 = _T_7871 ? 16'h40 : _T_8473; // @[Mux.scala 31:69:@4750.4]
  assign _T_8475 = _T_7868 ? 16'h20 : _T_8474; // @[Mux.scala 31:69:@4751.4]
  assign _T_8476 = _T_7865 ? 16'h10 : _T_8475; // @[Mux.scala 31:69:@4752.4]
  assign _T_8477 = _T_7862 ? 16'h8 : _T_8476; // @[Mux.scala 31:69:@4753.4]
  assign _T_8478 = _T_7859 ? 16'h4 : _T_8477; // @[Mux.scala 31:69:@4754.4]
  assign _T_8479 = _T_7856 ? 16'h2 : _T_8478; // @[Mux.scala 31:69:@4755.4]
  assign _T_8480 = _T_7853 ? 16'h1 : _T_8479; // @[Mux.scala 31:69:@4756.4]
  assign _T_8481 = _T_8480[0]; // @[OneHot.scala 66:30:@4757.4]
  assign _T_8482 = _T_8480[1]; // @[OneHot.scala 66:30:@4758.4]
  assign _T_8483 = _T_8480[2]; // @[OneHot.scala 66:30:@4759.4]
  assign _T_8484 = _T_8480[3]; // @[OneHot.scala 66:30:@4760.4]
  assign _T_8485 = _T_8480[4]; // @[OneHot.scala 66:30:@4761.4]
  assign _T_8486 = _T_8480[5]; // @[OneHot.scala 66:30:@4762.4]
  assign _T_8487 = _T_8480[6]; // @[OneHot.scala 66:30:@4763.4]
  assign _T_8488 = _T_8480[7]; // @[OneHot.scala 66:30:@4764.4]
  assign _T_8489 = _T_8480[8]; // @[OneHot.scala 66:30:@4765.4]
  assign _T_8490 = _T_8480[9]; // @[OneHot.scala 66:30:@4766.4]
  assign _T_8491 = _T_8480[10]; // @[OneHot.scala 66:30:@4767.4]
  assign _T_8492 = _T_8480[11]; // @[OneHot.scala 66:30:@4768.4]
  assign _T_8493 = _T_8480[12]; // @[OneHot.scala 66:30:@4769.4]
  assign _T_8494 = _T_8480[13]; // @[OneHot.scala 66:30:@4770.4]
  assign _T_8495 = _T_8480[14]; // @[OneHot.scala 66:30:@4771.4]
  assign _T_8496 = _T_8480[15]; // @[OneHot.scala 66:30:@4772.4]
  assign _T_8537 = _T_7853 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4790.4]
  assign _T_8538 = _T_7850 ? 16'h4000 : _T_8537; // @[Mux.scala 31:69:@4791.4]
  assign _T_8539 = _T_7847 ? 16'h2000 : _T_8538; // @[Mux.scala 31:69:@4792.4]
  assign _T_8540 = _T_7844 ? 16'h1000 : _T_8539; // @[Mux.scala 31:69:@4793.4]
  assign _T_8541 = _T_7841 ? 16'h800 : _T_8540; // @[Mux.scala 31:69:@4794.4]
  assign _T_8542 = _T_7838 ? 16'h400 : _T_8541; // @[Mux.scala 31:69:@4795.4]
  assign _T_8543 = _T_7835 ? 16'h200 : _T_8542; // @[Mux.scala 31:69:@4796.4]
  assign _T_8544 = _T_7880 ? 16'h100 : _T_8543; // @[Mux.scala 31:69:@4797.4]
  assign _T_8545 = _T_7877 ? 16'h80 : _T_8544; // @[Mux.scala 31:69:@4798.4]
  assign _T_8546 = _T_7874 ? 16'h40 : _T_8545; // @[Mux.scala 31:69:@4799.4]
  assign _T_8547 = _T_7871 ? 16'h20 : _T_8546; // @[Mux.scala 31:69:@4800.4]
  assign _T_8548 = _T_7868 ? 16'h10 : _T_8547; // @[Mux.scala 31:69:@4801.4]
  assign _T_8549 = _T_7865 ? 16'h8 : _T_8548; // @[Mux.scala 31:69:@4802.4]
  assign _T_8550 = _T_7862 ? 16'h4 : _T_8549; // @[Mux.scala 31:69:@4803.4]
  assign _T_8551 = _T_7859 ? 16'h2 : _T_8550; // @[Mux.scala 31:69:@4804.4]
  assign _T_8552 = _T_7856 ? 16'h1 : _T_8551; // @[Mux.scala 31:69:@4805.4]
  assign _T_8553 = _T_8552[0]; // @[OneHot.scala 66:30:@4806.4]
  assign _T_8554 = _T_8552[1]; // @[OneHot.scala 66:30:@4807.4]
  assign _T_8555 = _T_8552[2]; // @[OneHot.scala 66:30:@4808.4]
  assign _T_8556 = _T_8552[3]; // @[OneHot.scala 66:30:@4809.4]
  assign _T_8557 = _T_8552[4]; // @[OneHot.scala 66:30:@4810.4]
  assign _T_8558 = _T_8552[5]; // @[OneHot.scala 66:30:@4811.4]
  assign _T_8559 = _T_8552[6]; // @[OneHot.scala 66:30:@4812.4]
  assign _T_8560 = _T_8552[7]; // @[OneHot.scala 66:30:@4813.4]
  assign _T_8561 = _T_8552[8]; // @[OneHot.scala 66:30:@4814.4]
  assign _T_8562 = _T_8552[9]; // @[OneHot.scala 66:30:@4815.4]
  assign _T_8563 = _T_8552[10]; // @[OneHot.scala 66:30:@4816.4]
  assign _T_8564 = _T_8552[11]; // @[OneHot.scala 66:30:@4817.4]
  assign _T_8565 = _T_8552[12]; // @[OneHot.scala 66:30:@4818.4]
  assign _T_8566 = _T_8552[13]; // @[OneHot.scala 66:30:@4819.4]
  assign _T_8567 = _T_8552[14]; // @[OneHot.scala 66:30:@4820.4]
  assign _T_8568 = _T_8552[15]; // @[OneHot.scala 66:30:@4821.4]
  assign _T_8609 = _T_7856 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4839.4]
  assign _T_8610 = _T_7853 ? 16'h4000 : _T_8609; // @[Mux.scala 31:69:@4840.4]
  assign _T_8611 = _T_7850 ? 16'h2000 : _T_8610; // @[Mux.scala 31:69:@4841.4]
  assign _T_8612 = _T_7847 ? 16'h1000 : _T_8611; // @[Mux.scala 31:69:@4842.4]
  assign _T_8613 = _T_7844 ? 16'h800 : _T_8612; // @[Mux.scala 31:69:@4843.4]
  assign _T_8614 = _T_7841 ? 16'h400 : _T_8613; // @[Mux.scala 31:69:@4844.4]
  assign _T_8615 = _T_7838 ? 16'h200 : _T_8614; // @[Mux.scala 31:69:@4845.4]
  assign _T_8616 = _T_7835 ? 16'h100 : _T_8615; // @[Mux.scala 31:69:@4846.4]
  assign _T_8617 = _T_7880 ? 16'h80 : _T_8616; // @[Mux.scala 31:69:@4847.4]
  assign _T_8618 = _T_7877 ? 16'h40 : _T_8617; // @[Mux.scala 31:69:@4848.4]
  assign _T_8619 = _T_7874 ? 16'h20 : _T_8618; // @[Mux.scala 31:69:@4849.4]
  assign _T_8620 = _T_7871 ? 16'h10 : _T_8619; // @[Mux.scala 31:69:@4850.4]
  assign _T_8621 = _T_7868 ? 16'h8 : _T_8620; // @[Mux.scala 31:69:@4851.4]
  assign _T_8622 = _T_7865 ? 16'h4 : _T_8621; // @[Mux.scala 31:69:@4852.4]
  assign _T_8623 = _T_7862 ? 16'h2 : _T_8622; // @[Mux.scala 31:69:@4853.4]
  assign _T_8624 = _T_7859 ? 16'h1 : _T_8623; // @[Mux.scala 31:69:@4854.4]
  assign _T_8625 = _T_8624[0]; // @[OneHot.scala 66:30:@4855.4]
  assign _T_8626 = _T_8624[1]; // @[OneHot.scala 66:30:@4856.4]
  assign _T_8627 = _T_8624[2]; // @[OneHot.scala 66:30:@4857.4]
  assign _T_8628 = _T_8624[3]; // @[OneHot.scala 66:30:@4858.4]
  assign _T_8629 = _T_8624[4]; // @[OneHot.scala 66:30:@4859.4]
  assign _T_8630 = _T_8624[5]; // @[OneHot.scala 66:30:@4860.4]
  assign _T_8631 = _T_8624[6]; // @[OneHot.scala 66:30:@4861.4]
  assign _T_8632 = _T_8624[7]; // @[OneHot.scala 66:30:@4862.4]
  assign _T_8633 = _T_8624[8]; // @[OneHot.scala 66:30:@4863.4]
  assign _T_8634 = _T_8624[9]; // @[OneHot.scala 66:30:@4864.4]
  assign _T_8635 = _T_8624[10]; // @[OneHot.scala 66:30:@4865.4]
  assign _T_8636 = _T_8624[11]; // @[OneHot.scala 66:30:@4866.4]
  assign _T_8637 = _T_8624[12]; // @[OneHot.scala 66:30:@4867.4]
  assign _T_8638 = _T_8624[13]; // @[OneHot.scala 66:30:@4868.4]
  assign _T_8639 = _T_8624[14]; // @[OneHot.scala 66:30:@4869.4]
  assign _T_8640 = _T_8624[15]; // @[OneHot.scala 66:30:@4870.4]
  assign _T_8681 = _T_7859 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4888.4]
  assign _T_8682 = _T_7856 ? 16'h4000 : _T_8681; // @[Mux.scala 31:69:@4889.4]
  assign _T_8683 = _T_7853 ? 16'h2000 : _T_8682; // @[Mux.scala 31:69:@4890.4]
  assign _T_8684 = _T_7850 ? 16'h1000 : _T_8683; // @[Mux.scala 31:69:@4891.4]
  assign _T_8685 = _T_7847 ? 16'h800 : _T_8684; // @[Mux.scala 31:69:@4892.4]
  assign _T_8686 = _T_7844 ? 16'h400 : _T_8685; // @[Mux.scala 31:69:@4893.4]
  assign _T_8687 = _T_7841 ? 16'h200 : _T_8686; // @[Mux.scala 31:69:@4894.4]
  assign _T_8688 = _T_7838 ? 16'h100 : _T_8687; // @[Mux.scala 31:69:@4895.4]
  assign _T_8689 = _T_7835 ? 16'h80 : _T_8688; // @[Mux.scala 31:69:@4896.4]
  assign _T_8690 = _T_7880 ? 16'h40 : _T_8689; // @[Mux.scala 31:69:@4897.4]
  assign _T_8691 = _T_7877 ? 16'h20 : _T_8690; // @[Mux.scala 31:69:@4898.4]
  assign _T_8692 = _T_7874 ? 16'h10 : _T_8691; // @[Mux.scala 31:69:@4899.4]
  assign _T_8693 = _T_7871 ? 16'h8 : _T_8692; // @[Mux.scala 31:69:@4900.4]
  assign _T_8694 = _T_7868 ? 16'h4 : _T_8693; // @[Mux.scala 31:69:@4901.4]
  assign _T_8695 = _T_7865 ? 16'h2 : _T_8694; // @[Mux.scala 31:69:@4902.4]
  assign _T_8696 = _T_7862 ? 16'h1 : _T_8695; // @[Mux.scala 31:69:@4903.4]
  assign _T_8697 = _T_8696[0]; // @[OneHot.scala 66:30:@4904.4]
  assign _T_8698 = _T_8696[1]; // @[OneHot.scala 66:30:@4905.4]
  assign _T_8699 = _T_8696[2]; // @[OneHot.scala 66:30:@4906.4]
  assign _T_8700 = _T_8696[3]; // @[OneHot.scala 66:30:@4907.4]
  assign _T_8701 = _T_8696[4]; // @[OneHot.scala 66:30:@4908.4]
  assign _T_8702 = _T_8696[5]; // @[OneHot.scala 66:30:@4909.4]
  assign _T_8703 = _T_8696[6]; // @[OneHot.scala 66:30:@4910.4]
  assign _T_8704 = _T_8696[7]; // @[OneHot.scala 66:30:@4911.4]
  assign _T_8705 = _T_8696[8]; // @[OneHot.scala 66:30:@4912.4]
  assign _T_8706 = _T_8696[9]; // @[OneHot.scala 66:30:@4913.4]
  assign _T_8707 = _T_8696[10]; // @[OneHot.scala 66:30:@4914.4]
  assign _T_8708 = _T_8696[11]; // @[OneHot.scala 66:30:@4915.4]
  assign _T_8709 = _T_8696[12]; // @[OneHot.scala 66:30:@4916.4]
  assign _T_8710 = _T_8696[13]; // @[OneHot.scala 66:30:@4917.4]
  assign _T_8711 = _T_8696[14]; // @[OneHot.scala 66:30:@4918.4]
  assign _T_8712 = _T_8696[15]; // @[OneHot.scala 66:30:@4919.4]
  assign _T_8753 = _T_7862 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4937.4]
  assign _T_8754 = _T_7859 ? 16'h4000 : _T_8753; // @[Mux.scala 31:69:@4938.4]
  assign _T_8755 = _T_7856 ? 16'h2000 : _T_8754; // @[Mux.scala 31:69:@4939.4]
  assign _T_8756 = _T_7853 ? 16'h1000 : _T_8755; // @[Mux.scala 31:69:@4940.4]
  assign _T_8757 = _T_7850 ? 16'h800 : _T_8756; // @[Mux.scala 31:69:@4941.4]
  assign _T_8758 = _T_7847 ? 16'h400 : _T_8757; // @[Mux.scala 31:69:@4942.4]
  assign _T_8759 = _T_7844 ? 16'h200 : _T_8758; // @[Mux.scala 31:69:@4943.4]
  assign _T_8760 = _T_7841 ? 16'h100 : _T_8759; // @[Mux.scala 31:69:@4944.4]
  assign _T_8761 = _T_7838 ? 16'h80 : _T_8760; // @[Mux.scala 31:69:@4945.4]
  assign _T_8762 = _T_7835 ? 16'h40 : _T_8761; // @[Mux.scala 31:69:@4946.4]
  assign _T_8763 = _T_7880 ? 16'h20 : _T_8762; // @[Mux.scala 31:69:@4947.4]
  assign _T_8764 = _T_7877 ? 16'h10 : _T_8763; // @[Mux.scala 31:69:@4948.4]
  assign _T_8765 = _T_7874 ? 16'h8 : _T_8764; // @[Mux.scala 31:69:@4949.4]
  assign _T_8766 = _T_7871 ? 16'h4 : _T_8765; // @[Mux.scala 31:69:@4950.4]
  assign _T_8767 = _T_7868 ? 16'h2 : _T_8766; // @[Mux.scala 31:69:@4951.4]
  assign _T_8768 = _T_7865 ? 16'h1 : _T_8767; // @[Mux.scala 31:69:@4952.4]
  assign _T_8769 = _T_8768[0]; // @[OneHot.scala 66:30:@4953.4]
  assign _T_8770 = _T_8768[1]; // @[OneHot.scala 66:30:@4954.4]
  assign _T_8771 = _T_8768[2]; // @[OneHot.scala 66:30:@4955.4]
  assign _T_8772 = _T_8768[3]; // @[OneHot.scala 66:30:@4956.4]
  assign _T_8773 = _T_8768[4]; // @[OneHot.scala 66:30:@4957.4]
  assign _T_8774 = _T_8768[5]; // @[OneHot.scala 66:30:@4958.4]
  assign _T_8775 = _T_8768[6]; // @[OneHot.scala 66:30:@4959.4]
  assign _T_8776 = _T_8768[7]; // @[OneHot.scala 66:30:@4960.4]
  assign _T_8777 = _T_8768[8]; // @[OneHot.scala 66:30:@4961.4]
  assign _T_8778 = _T_8768[9]; // @[OneHot.scala 66:30:@4962.4]
  assign _T_8779 = _T_8768[10]; // @[OneHot.scala 66:30:@4963.4]
  assign _T_8780 = _T_8768[11]; // @[OneHot.scala 66:30:@4964.4]
  assign _T_8781 = _T_8768[12]; // @[OneHot.scala 66:30:@4965.4]
  assign _T_8782 = _T_8768[13]; // @[OneHot.scala 66:30:@4966.4]
  assign _T_8783 = _T_8768[14]; // @[OneHot.scala 66:30:@4967.4]
  assign _T_8784 = _T_8768[15]; // @[OneHot.scala 66:30:@4968.4]
  assign _T_8825 = _T_7865 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@4986.4]
  assign _T_8826 = _T_7862 ? 16'h4000 : _T_8825; // @[Mux.scala 31:69:@4987.4]
  assign _T_8827 = _T_7859 ? 16'h2000 : _T_8826; // @[Mux.scala 31:69:@4988.4]
  assign _T_8828 = _T_7856 ? 16'h1000 : _T_8827; // @[Mux.scala 31:69:@4989.4]
  assign _T_8829 = _T_7853 ? 16'h800 : _T_8828; // @[Mux.scala 31:69:@4990.4]
  assign _T_8830 = _T_7850 ? 16'h400 : _T_8829; // @[Mux.scala 31:69:@4991.4]
  assign _T_8831 = _T_7847 ? 16'h200 : _T_8830; // @[Mux.scala 31:69:@4992.4]
  assign _T_8832 = _T_7844 ? 16'h100 : _T_8831; // @[Mux.scala 31:69:@4993.4]
  assign _T_8833 = _T_7841 ? 16'h80 : _T_8832; // @[Mux.scala 31:69:@4994.4]
  assign _T_8834 = _T_7838 ? 16'h40 : _T_8833; // @[Mux.scala 31:69:@4995.4]
  assign _T_8835 = _T_7835 ? 16'h20 : _T_8834; // @[Mux.scala 31:69:@4996.4]
  assign _T_8836 = _T_7880 ? 16'h10 : _T_8835; // @[Mux.scala 31:69:@4997.4]
  assign _T_8837 = _T_7877 ? 16'h8 : _T_8836; // @[Mux.scala 31:69:@4998.4]
  assign _T_8838 = _T_7874 ? 16'h4 : _T_8837; // @[Mux.scala 31:69:@4999.4]
  assign _T_8839 = _T_7871 ? 16'h2 : _T_8838; // @[Mux.scala 31:69:@5000.4]
  assign _T_8840 = _T_7868 ? 16'h1 : _T_8839; // @[Mux.scala 31:69:@5001.4]
  assign _T_8841 = _T_8840[0]; // @[OneHot.scala 66:30:@5002.4]
  assign _T_8842 = _T_8840[1]; // @[OneHot.scala 66:30:@5003.4]
  assign _T_8843 = _T_8840[2]; // @[OneHot.scala 66:30:@5004.4]
  assign _T_8844 = _T_8840[3]; // @[OneHot.scala 66:30:@5005.4]
  assign _T_8845 = _T_8840[4]; // @[OneHot.scala 66:30:@5006.4]
  assign _T_8846 = _T_8840[5]; // @[OneHot.scala 66:30:@5007.4]
  assign _T_8847 = _T_8840[6]; // @[OneHot.scala 66:30:@5008.4]
  assign _T_8848 = _T_8840[7]; // @[OneHot.scala 66:30:@5009.4]
  assign _T_8849 = _T_8840[8]; // @[OneHot.scala 66:30:@5010.4]
  assign _T_8850 = _T_8840[9]; // @[OneHot.scala 66:30:@5011.4]
  assign _T_8851 = _T_8840[10]; // @[OneHot.scala 66:30:@5012.4]
  assign _T_8852 = _T_8840[11]; // @[OneHot.scala 66:30:@5013.4]
  assign _T_8853 = _T_8840[12]; // @[OneHot.scala 66:30:@5014.4]
  assign _T_8854 = _T_8840[13]; // @[OneHot.scala 66:30:@5015.4]
  assign _T_8855 = _T_8840[14]; // @[OneHot.scala 66:30:@5016.4]
  assign _T_8856 = _T_8840[15]; // @[OneHot.scala 66:30:@5017.4]
  assign _T_8897 = _T_7868 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5035.4]
  assign _T_8898 = _T_7865 ? 16'h4000 : _T_8897; // @[Mux.scala 31:69:@5036.4]
  assign _T_8899 = _T_7862 ? 16'h2000 : _T_8898; // @[Mux.scala 31:69:@5037.4]
  assign _T_8900 = _T_7859 ? 16'h1000 : _T_8899; // @[Mux.scala 31:69:@5038.4]
  assign _T_8901 = _T_7856 ? 16'h800 : _T_8900; // @[Mux.scala 31:69:@5039.4]
  assign _T_8902 = _T_7853 ? 16'h400 : _T_8901; // @[Mux.scala 31:69:@5040.4]
  assign _T_8903 = _T_7850 ? 16'h200 : _T_8902; // @[Mux.scala 31:69:@5041.4]
  assign _T_8904 = _T_7847 ? 16'h100 : _T_8903; // @[Mux.scala 31:69:@5042.4]
  assign _T_8905 = _T_7844 ? 16'h80 : _T_8904; // @[Mux.scala 31:69:@5043.4]
  assign _T_8906 = _T_7841 ? 16'h40 : _T_8905; // @[Mux.scala 31:69:@5044.4]
  assign _T_8907 = _T_7838 ? 16'h20 : _T_8906; // @[Mux.scala 31:69:@5045.4]
  assign _T_8908 = _T_7835 ? 16'h10 : _T_8907; // @[Mux.scala 31:69:@5046.4]
  assign _T_8909 = _T_7880 ? 16'h8 : _T_8908; // @[Mux.scala 31:69:@5047.4]
  assign _T_8910 = _T_7877 ? 16'h4 : _T_8909; // @[Mux.scala 31:69:@5048.4]
  assign _T_8911 = _T_7874 ? 16'h2 : _T_8910; // @[Mux.scala 31:69:@5049.4]
  assign _T_8912 = _T_7871 ? 16'h1 : _T_8911; // @[Mux.scala 31:69:@5050.4]
  assign _T_8913 = _T_8912[0]; // @[OneHot.scala 66:30:@5051.4]
  assign _T_8914 = _T_8912[1]; // @[OneHot.scala 66:30:@5052.4]
  assign _T_8915 = _T_8912[2]; // @[OneHot.scala 66:30:@5053.4]
  assign _T_8916 = _T_8912[3]; // @[OneHot.scala 66:30:@5054.4]
  assign _T_8917 = _T_8912[4]; // @[OneHot.scala 66:30:@5055.4]
  assign _T_8918 = _T_8912[5]; // @[OneHot.scala 66:30:@5056.4]
  assign _T_8919 = _T_8912[6]; // @[OneHot.scala 66:30:@5057.4]
  assign _T_8920 = _T_8912[7]; // @[OneHot.scala 66:30:@5058.4]
  assign _T_8921 = _T_8912[8]; // @[OneHot.scala 66:30:@5059.4]
  assign _T_8922 = _T_8912[9]; // @[OneHot.scala 66:30:@5060.4]
  assign _T_8923 = _T_8912[10]; // @[OneHot.scala 66:30:@5061.4]
  assign _T_8924 = _T_8912[11]; // @[OneHot.scala 66:30:@5062.4]
  assign _T_8925 = _T_8912[12]; // @[OneHot.scala 66:30:@5063.4]
  assign _T_8926 = _T_8912[13]; // @[OneHot.scala 66:30:@5064.4]
  assign _T_8927 = _T_8912[14]; // @[OneHot.scala 66:30:@5065.4]
  assign _T_8928 = _T_8912[15]; // @[OneHot.scala 66:30:@5066.4]
  assign _T_8969 = _T_7871 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5084.4]
  assign _T_8970 = _T_7868 ? 16'h4000 : _T_8969; // @[Mux.scala 31:69:@5085.4]
  assign _T_8971 = _T_7865 ? 16'h2000 : _T_8970; // @[Mux.scala 31:69:@5086.4]
  assign _T_8972 = _T_7862 ? 16'h1000 : _T_8971; // @[Mux.scala 31:69:@5087.4]
  assign _T_8973 = _T_7859 ? 16'h800 : _T_8972; // @[Mux.scala 31:69:@5088.4]
  assign _T_8974 = _T_7856 ? 16'h400 : _T_8973; // @[Mux.scala 31:69:@5089.4]
  assign _T_8975 = _T_7853 ? 16'h200 : _T_8974; // @[Mux.scala 31:69:@5090.4]
  assign _T_8976 = _T_7850 ? 16'h100 : _T_8975; // @[Mux.scala 31:69:@5091.4]
  assign _T_8977 = _T_7847 ? 16'h80 : _T_8976; // @[Mux.scala 31:69:@5092.4]
  assign _T_8978 = _T_7844 ? 16'h40 : _T_8977; // @[Mux.scala 31:69:@5093.4]
  assign _T_8979 = _T_7841 ? 16'h20 : _T_8978; // @[Mux.scala 31:69:@5094.4]
  assign _T_8980 = _T_7838 ? 16'h10 : _T_8979; // @[Mux.scala 31:69:@5095.4]
  assign _T_8981 = _T_7835 ? 16'h8 : _T_8980; // @[Mux.scala 31:69:@5096.4]
  assign _T_8982 = _T_7880 ? 16'h4 : _T_8981; // @[Mux.scala 31:69:@5097.4]
  assign _T_8983 = _T_7877 ? 16'h2 : _T_8982; // @[Mux.scala 31:69:@5098.4]
  assign _T_8984 = _T_7874 ? 16'h1 : _T_8983; // @[Mux.scala 31:69:@5099.4]
  assign _T_8985 = _T_8984[0]; // @[OneHot.scala 66:30:@5100.4]
  assign _T_8986 = _T_8984[1]; // @[OneHot.scala 66:30:@5101.4]
  assign _T_8987 = _T_8984[2]; // @[OneHot.scala 66:30:@5102.4]
  assign _T_8988 = _T_8984[3]; // @[OneHot.scala 66:30:@5103.4]
  assign _T_8989 = _T_8984[4]; // @[OneHot.scala 66:30:@5104.4]
  assign _T_8990 = _T_8984[5]; // @[OneHot.scala 66:30:@5105.4]
  assign _T_8991 = _T_8984[6]; // @[OneHot.scala 66:30:@5106.4]
  assign _T_8992 = _T_8984[7]; // @[OneHot.scala 66:30:@5107.4]
  assign _T_8993 = _T_8984[8]; // @[OneHot.scala 66:30:@5108.4]
  assign _T_8994 = _T_8984[9]; // @[OneHot.scala 66:30:@5109.4]
  assign _T_8995 = _T_8984[10]; // @[OneHot.scala 66:30:@5110.4]
  assign _T_8996 = _T_8984[11]; // @[OneHot.scala 66:30:@5111.4]
  assign _T_8997 = _T_8984[12]; // @[OneHot.scala 66:30:@5112.4]
  assign _T_8998 = _T_8984[13]; // @[OneHot.scala 66:30:@5113.4]
  assign _T_8999 = _T_8984[14]; // @[OneHot.scala 66:30:@5114.4]
  assign _T_9000 = _T_8984[15]; // @[OneHot.scala 66:30:@5115.4]
  assign _T_9041 = _T_7874 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5133.4]
  assign _T_9042 = _T_7871 ? 16'h4000 : _T_9041; // @[Mux.scala 31:69:@5134.4]
  assign _T_9043 = _T_7868 ? 16'h2000 : _T_9042; // @[Mux.scala 31:69:@5135.4]
  assign _T_9044 = _T_7865 ? 16'h1000 : _T_9043; // @[Mux.scala 31:69:@5136.4]
  assign _T_9045 = _T_7862 ? 16'h800 : _T_9044; // @[Mux.scala 31:69:@5137.4]
  assign _T_9046 = _T_7859 ? 16'h400 : _T_9045; // @[Mux.scala 31:69:@5138.4]
  assign _T_9047 = _T_7856 ? 16'h200 : _T_9046; // @[Mux.scala 31:69:@5139.4]
  assign _T_9048 = _T_7853 ? 16'h100 : _T_9047; // @[Mux.scala 31:69:@5140.4]
  assign _T_9049 = _T_7850 ? 16'h80 : _T_9048; // @[Mux.scala 31:69:@5141.4]
  assign _T_9050 = _T_7847 ? 16'h40 : _T_9049; // @[Mux.scala 31:69:@5142.4]
  assign _T_9051 = _T_7844 ? 16'h20 : _T_9050; // @[Mux.scala 31:69:@5143.4]
  assign _T_9052 = _T_7841 ? 16'h10 : _T_9051; // @[Mux.scala 31:69:@5144.4]
  assign _T_9053 = _T_7838 ? 16'h8 : _T_9052; // @[Mux.scala 31:69:@5145.4]
  assign _T_9054 = _T_7835 ? 16'h4 : _T_9053; // @[Mux.scala 31:69:@5146.4]
  assign _T_9055 = _T_7880 ? 16'h2 : _T_9054; // @[Mux.scala 31:69:@5147.4]
  assign _T_9056 = _T_7877 ? 16'h1 : _T_9055; // @[Mux.scala 31:69:@5148.4]
  assign _T_9057 = _T_9056[0]; // @[OneHot.scala 66:30:@5149.4]
  assign _T_9058 = _T_9056[1]; // @[OneHot.scala 66:30:@5150.4]
  assign _T_9059 = _T_9056[2]; // @[OneHot.scala 66:30:@5151.4]
  assign _T_9060 = _T_9056[3]; // @[OneHot.scala 66:30:@5152.4]
  assign _T_9061 = _T_9056[4]; // @[OneHot.scala 66:30:@5153.4]
  assign _T_9062 = _T_9056[5]; // @[OneHot.scala 66:30:@5154.4]
  assign _T_9063 = _T_9056[6]; // @[OneHot.scala 66:30:@5155.4]
  assign _T_9064 = _T_9056[7]; // @[OneHot.scala 66:30:@5156.4]
  assign _T_9065 = _T_9056[8]; // @[OneHot.scala 66:30:@5157.4]
  assign _T_9066 = _T_9056[9]; // @[OneHot.scala 66:30:@5158.4]
  assign _T_9067 = _T_9056[10]; // @[OneHot.scala 66:30:@5159.4]
  assign _T_9068 = _T_9056[11]; // @[OneHot.scala 66:30:@5160.4]
  assign _T_9069 = _T_9056[12]; // @[OneHot.scala 66:30:@5161.4]
  assign _T_9070 = _T_9056[13]; // @[OneHot.scala 66:30:@5162.4]
  assign _T_9071 = _T_9056[14]; // @[OneHot.scala 66:30:@5163.4]
  assign _T_9072 = _T_9056[15]; // @[OneHot.scala 66:30:@5164.4]
  assign _T_9113 = _T_7877 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5182.4]
  assign _T_9114 = _T_7874 ? 16'h4000 : _T_9113; // @[Mux.scala 31:69:@5183.4]
  assign _T_9115 = _T_7871 ? 16'h2000 : _T_9114; // @[Mux.scala 31:69:@5184.4]
  assign _T_9116 = _T_7868 ? 16'h1000 : _T_9115; // @[Mux.scala 31:69:@5185.4]
  assign _T_9117 = _T_7865 ? 16'h800 : _T_9116; // @[Mux.scala 31:69:@5186.4]
  assign _T_9118 = _T_7862 ? 16'h400 : _T_9117; // @[Mux.scala 31:69:@5187.4]
  assign _T_9119 = _T_7859 ? 16'h200 : _T_9118; // @[Mux.scala 31:69:@5188.4]
  assign _T_9120 = _T_7856 ? 16'h100 : _T_9119; // @[Mux.scala 31:69:@5189.4]
  assign _T_9121 = _T_7853 ? 16'h80 : _T_9120; // @[Mux.scala 31:69:@5190.4]
  assign _T_9122 = _T_7850 ? 16'h40 : _T_9121; // @[Mux.scala 31:69:@5191.4]
  assign _T_9123 = _T_7847 ? 16'h20 : _T_9122; // @[Mux.scala 31:69:@5192.4]
  assign _T_9124 = _T_7844 ? 16'h10 : _T_9123; // @[Mux.scala 31:69:@5193.4]
  assign _T_9125 = _T_7841 ? 16'h8 : _T_9124; // @[Mux.scala 31:69:@5194.4]
  assign _T_9126 = _T_7838 ? 16'h4 : _T_9125; // @[Mux.scala 31:69:@5195.4]
  assign _T_9127 = _T_7835 ? 16'h2 : _T_9126; // @[Mux.scala 31:69:@5196.4]
  assign _T_9128 = _T_7880 ? 16'h1 : _T_9127; // @[Mux.scala 31:69:@5197.4]
  assign _T_9129 = _T_9128[0]; // @[OneHot.scala 66:30:@5198.4]
  assign _T_9130 = _T_9128[1]; // @[OneHot.scala 66:30:@5199.4]
  assign _T_9131 = _T_9128[2]; // @[OneHot.scala 66:30:@5200.4]
  assign _T_9132 = _T_9128[3]; // @[OneHot.scala 66:30:@5201.4]
  assign _T_9133 = _T_9128[4]; // @[OneHot.scala 66:30:@5202.4]
  assign _T_9134 = _T_9128[5]; // @[OneHot.scala 66:30:@5203.4]
  assign _T_9135 = _T_9128[6]; // @[OneHot.scala 66:30:@5204.4]
  assign _T_9136 = _T_9128[7]; // @[OneHot.scala 66:30:@5205.4]
  assign _T_9137 = _T_9128[8]; // @[OneHot.scala 66:30:@5206.4]
  assign _T_9138 = _T_9128[9]; // @[OneHot.scala 66:30:@5207.4]
  assign _T_9139 = _T_9128[10]; // @[OneHot.scala 66:30:@5208.4]
  assign _T_9140 = _T_9128[11]; // @[OneHot.scala 66:30:@5209.4]
  assign _T_9141 = _T_9128[12]; // @[OneHot.scala 66:30:@5210.4]
  assign _T_9142 = _T_9128[13]; // @[OneHot.scala 66:30:@5211.4]
  assign _T_9143 = _T_9128[14]; // @[OneHot.scala 66:30:@5212.4]
  assign _T_9144 = _T_9128[15]; // @[OneHot.scala 66:30:@5213.4]
  assign _T_9209 = {_T_8056,_T_8055,_T_8054,_T_8053,_T_8052,_T_8051,_T_8050,_T_8049}; // @[Mux.scala 19:72:@5237.4]
  assign _T_9217 = {_T_8064,_T_8063,_T_8062,_T_8061,_T_8060,_T_8059,_T_8058,_T_8057,_T_9209}; // @[Mux.scala 19:72:@5245.4]
  assign _T_9219 = _T_4521 ? _T_9217 : 16'h0; // @[Mux.scala 19:72:@5246.4]
  assign _T_9226 = {_T_8127,_T_8126,_T_8125,_T_8124,_T_8123,_T_8122,_T_8121,_T_8136}; // @[Mux.scala 19:72:@5253.4]
  assign _T_9234 = {_T_8135,_T_8134,_T_8133,_T_8132,_T_8131,_T_8130,_T_8129,_T_8128,_T_9226}; // @[Mux.scala 19:72:@5261.4]
  assign _T_9236 = _T_4522 ? _T_9234 : 16'h0; // @[Mux.scala 19:72:@5262.4]
  assign _T_9243 = {_T_8198,_T_8197,_T_8196,_T_8195,_T_8194,_T_8193,_T_8208,_T_8207}; // @[Mux.scala 19:72:@5269.4]
  assign _T_9251 = {_T_8206,_T_8205,_T_8204,_T_8203,_T_8202,_T_8201,_T_8200,_T_8199,_T_9243}; // @[Mux.scala 19:72:@5277.4]
  assign _T_9253 = _T_4523 ? _T_9251 : 16'h0; // @[Mux.scala 19:72:@5278.4]
  assign _T_9260 = {_T_8269,_T_8268,_T_8267,_T_8266,_T_8265,_T_8280,_T_8279,_T_8278}; // @[Mux.scala 19:72:@5285.4]
  assign _T_9268 = {_T_8277,_T_8276,_T_8275,_T_8274,_T_8273,_T_8272,_T_8271,_T_8270,_T_9260}; // @[Mux.scala 19:72:@5293.4]
  assign _T_9270 = _T_4524 ? _T_9268 : 16'h0; // @[Mux.scala 19:72:@5294.4]
  assign _T_9277 = {_T_8340,_T_8339,_T_8338,_T_8337,_T_8352,_T_8351,_T_8350,_T_8349}; // @[Mux.scala 19:72:@5301.4]
  assign _T_9285 = {_T_8348,_T_8347,_T_8346,_T_8345,_T_8344,_T_8343,_T_8342,_T_8341,_T_9277}; // @[Mux.scala 19:72:@5309.4]
  assign _T_9287 = _T_4525 ? _T_9285 : 16'h0; // @[Mux.scala 19:72:@5310.4]
  assign _T_9294 = {_T_8411,_T_8410,_T_8409,_T_8424,_T_8423,_T_8422,_T_8421,_T_8420}; // @[Mux.scala 19:72:@5317.4]
  assign _T_9302 = {_T_8419,_T_8418,_T_8417,_T_8416,_T_8415,_T_8414,_T_8413,_T_8412,_T_9294}; // @[Mux.scala 19:72:@5325.4]
  assign _T_9304 = _T_4526 ? _T_9302 : 16'h0; // @[Mux.scala 19:72:@5326.4]
  assign _T_9311 = {_T_8482,_T_8481,_T_8496,_T_8495,_T_8494,_T_8493,_T_8492,_T_8491}; // @[Mux.scala 19:72:@5333.4]
  assign _T_9319 = {_T_8490,_T_8489,_T_8488,_T_8487,_T_8486,_T_8485,_T_8484,_T_8483,_T_9311}; // @[Mux.scala 19:72:@5341.4]
  assign _T_9321 = _T_4527 ? _T_9319 : 16'h0; // @[Mux.scala 19:72:@5342.4]
  assign _T_9328 = {_T_8553,_T_8568,_T_8567,_T_8566,_T_8565,_T_8564,_T_8563,_T_8562}; // @[Mux.scala 19:72:@5349.4]
  assign _T_9336 = {_T_8561,_T_8560,_T_8559,_T_8558,_T_8557,_T_8556,_T_8555,_T_8554,_T_9328}; // @[Mux.scala 19:72:@5357.4]
  assign _T_9338 = _T_4528 ? _T_9336 : 16'h0; // @[Mux.scala 19:72:@5358.4]
  assign _T_9345 = {_T_8640,_T_8639,_T_8638,_T_8637,_T_8636,_T_8635,_T_8634,_T_8633}; // @[Mux.scala 19:72:@5365.4]
  assign _T_9353 = {_T_8632,_T_8631,_T_8630,_T_8629,_T_8628,_T_8627,_T_8626,_T_8625,_T_9345}; // @[Mux.scala 19:72:@5373.4]
  assign _T_9355 = _T_4529 ? _T_9353 : 16'h0; // @[Mux.scala 19:72:@5374.4]
  assign _T_9362 = {_T_8711,_T_8710,_T_8709,_T_8708,_T_8707,_T_8706,_T_8705,_T_8704}; // @[Mux.scala 19:72:@5381.4]
  assign _T_9370 = {_T_8703,_T_8702,_T_8701,_T_8700,_T_8699,_T_8698,_T_8697,_T_8712,_T_9362}; // @[Mux.scala 19:72:@5389.4]
  assign _T_9372 = _T_4530 ? _T_9370 : 16'h0; // @[Mux.scala 19:72:@5390.4]
  assign _T_9379 = {_T_8782,_T_8781,_T_8780,_T_8779,_T_8778,_T_8777,_T_8776,_T_8775}; // @[Mux.scala 19:72:@5397.4]
  assign _T_9387 = {_T_8774,_T_8773,_T_8772,_T_8771,_T_8770,_T_8769,_T_8784,_T_8783,_T_9379}; // @[Mux.scala 19:72:@5405.4]
  assign _T_9389 = _T_4531 ? _T_9387 : 16'h0; // @[Mux.scala 19:72:@5406.4]
  assign _T_9396 = {_T_8853,_T_8852,_T_8851,_T_8850,_T_8849,_T_8848,_T_8847,_T_8846}; // @[Mux.scala 19:72:@5413.4]
  assign _T_9404 = {_T_8845,_T_8844,_T_8843,_T_8842,_T_8841,_T_8856,_T_8855,_T_8854,_T_9396}; // @[Mux.scala 19:72:@5421.4]
  assign _T_9406 = _T_4532 ? _T_9404 : 16'h0; // @[Mux.scala 19:72:@5422.4]
  assign _T_9413 = {_T_8924,_T_8923,_T_8922,_T_8921,_T_8920,_T_8919,_T_8918,_T_8917}; // @[Mux.scala 19:72:@5429.4]
  assign _T_9421 = {_T_8916,_T_8915,_T_8914,_T_8913,_T_8928,_T_8927,_T_8926,_T_8925,_T_9413}; // @[Mux.scala 19:72:@5437.4]
  assign _T_9423 = _T_4533 ? _T_9421 : 16'h0; // @[Mux.scala 19:72:@5438.4]
  assign _T_9430 = {_T_8995,_T_8994,_T_8993,_T_8992,_T_8991,_T_8990,_T_8989,_T_8988}; // @[Mux.scala 19:72:@5445.4]
  assign _T_9438 = {_T_8987,_T_8986,_T_8985,_T_9000,_T_8999,_T_8998,_T_8997,_T_8996,_T_9430}; // @[Mux.scala 19:72:@5453.4]
  assign _T_9440 = _T_4534 ? _T_9438 : 16'h0; // @[Mux.scala 19:72:@5454.4]
  assign _T_9447 = {_T_9066,_T_9065,_T_9064,_T_9063,_T_9062,_T_9061,_T_9060,_T_9059}; // @[Mux.scala 19:72:@5461.4]
  assign _T_9455 = {_T_9058,_T_9057,_T_9072,_T_9071,_T_9070,_T_9069,_T_9068,_T_9067,_T_9447}; // @[Mux.scala 19:72:@5469.4]
  assign _T_9457 = _T_4535 ? _T_9455 : 16'h0; // @[Mux.scala 19:72:@5470.4]
  assign _T_9464 = {_T_9137,_T_9136,_T_9135,_T_9134,_T_9133,_T_9132,_T_9131,_T_9130}; // @[Mux.scala 19:72:@5477.4]
  assign _T_9472 = {_T_9129,_T_9144,_T_9143,_T_9142,_T_9141,_T_9140,_T_9139,_T_9138,_T_9464}; // @[Mux.scala 19:72:@5485.4]
  assign _T_9474 = _T_4536 ? _T_9472 : 16'h0; // @[Mux.scala 19:72:@5486.4]
  assign _T_9475 = _T_9219 | _T_9236; // @[Mux.scala 19:72:@5487.4]
  assign _T_9476 = _T_9475 | _T_9253; // @[Mux.scala 19:72:@5488.4]
  assign _T_9477 = _T_9476 | _T_9270; // @[Mux.scala 19:72:@5489.4]
  assign _T_9478 = _T_9477 | _T_9287; // @[Mux.scala 19:72:@5490.4]
  assign _T_9479 = _T_9478 | _T_9304; // @[Mux.scala 19:72:@5491.4]
  assign _T_9480 = _T_9479 | _T_9321; // @[Mux.scala 19:72:@5492.4]
  assign _T_9481 = _T_9480 | _T_9338; // @[Mux.scala 19:72:@5493.4]
  assign _T_9482 = _T_9481 | _T_9355; // @[Mux.scala 19:72:@5494.4]
  assign _T_9483 = _T_9482 | _T_9372; // @[Mux.scala 19:72:@5495.4]
  assign _T_9484 = _T_9483 | _T_9389; // @[Mux.scala 19:72:@5496.4]
  assign _T_9485 = _T_9484 | _T_9406; // @[Mux.scala 19:72:@5497.4]
  assign _T_9486 = _T_9485 | _T_9423; // @[Mux.scala 19:72:@5498.4]
  assign _T_9487 = _T_9486 | _T_9440; // @[Mux.scala 19:72:@5499.4]
  assign _T_9488 = _T_9487 | _T_9457; // @[Mux.scala 19:72:@5500.4]
  assign _T_9489 = _T_9488 | _T_9474; // @[Mux.scala 19:72:@5501.4]
  assign inputAddrPriorityPorts_1_0 = _T_9489[0]; // @[Mux.scala 19:72:@5505.4]
  assign inputAddrPriorityPorts_1_1 = _T_9489[1]; // @[Mux.scala 19:72:@5507.4]
  assign inputAddrPriorityPorts_1_2 = _T_9489[2]; // @[Mux.scala 19:72:@5509.4]
  assign inputAddrPriorityPorts_1_3 = _T_9489[3]; // @[Mux.scala 19:72:@5511.4]
  assign inputAddrPriorityPorts_1_4 = _T_9489[4]; // @[Mux.scala 19:72:@5513.4]
  assign inputAddrPriorityPorts_1_5 = _T_9489[5]; // @[Mux.scala 19:72:@5515.4]
  assign inputAddrPriorityPorts_1_6 = _T_9489[6]; // @[Mux.scala 19:72:@5517.4]
  assign inputAddrPriorityPorts_1_7 = _T_9489[7]; // @[Mux.scala 19:72:@5519.4]
  assign inputAddrPriorityPorts_1_8 = _T_9489[8]; // @[Mux.scala 19:72:@5521.4]
  assign inputAddrPriorityPorts_1_9 = _T_9489[9]; // @[Mux.scala 19:72:@5523.4]
  assign inputAddrPriorityPorts_1_10 = _T_9489[10]; // @[Mux.scala 19:72:@5525.4]
  assign inputAddrPriorityPorts_1_11 = _T_9489[11]; // @[Mux.scala 19:72:@5527.4]
  assign inputAddrPriorityPorts_1_12 = _T_9489[12]; // @[Mux.scala 19:72:@5529.4]
  assign inputAddrPriorityPorts_1_13 = _T_9489[13]; // @[Mux.scala 19:72:@5531.4]
  assign inputAddrPriorityPorts_1_14 = _T_9489[14]; // @[Mux.scala 19:72:@5533.4]
  assign inputAddrPriorityPorts_1_15 = _T_9489[15]; // @[Mux.scala 19:72:@5535.4]
  assign _T_9691 = _T_7950 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5589.4]
  assign _T_9692 = _T_7947 ? 16'h4000 : _T_9691; // @[Mux.scala 31:69:@5590.4]
  assign _T_9693 = _T_7944 ? 16'h2000 : _T_9692; // @[Mux.scala 31:69:@5591.4]
  assign _T_9694 = _T_7941 ? 16'h1000 : _T_9693; // @[Mux.scala 31:69:@5592.4]
  assign _T_9695 = _T_7938 ? 16'h800 : _T_9694; // @[Mux.scala 31:69:@5593.4]
  assign _T_9696 = _T_7935 ? 16'h400 : _T_9695; // @[Mux.scala 31:69:@5594.4]
  assign _T_9697 = _T_7932 ? 16'h200 : _T_9696; // @[Mux.scala 31:69:@5595.4]
  assign _T_9698 = _T_7929 ? 16'h100 : _T_9697; // @[Mux.scala 31:69:@5596.4]
  assign _T_9699 = _T_7926 ? 16'h80 : _T_9698; // @[Mux.scala 31:69:@5597.4]
  assign _T_9700 = _T_7923 ? 16'h40 : _T_9699; // @[Mux.scala 31:69:@5598.4]
  assign _T_9701 = _T_7920 ? 16'h20 : _T_9700; // @[Mux.scala 31:69:@5599.4]
  assign _T_9702 = _T_7917 ? 16'h10 : _T_9701; // @[Mux.scala 31:69:@5600.4]
  assign _T_9703 = _T_7914 ? 16'h8 : _T_9702; // @[Mux.scala 31:69:@5601.4]
  assign _T_9704 = _T_7911 ? 16'h4 : _T_9703; // @[Mux.scala 31:69:@5602.4]
  assign _T_9705 = _T_7908 ? 16'h2 : _T_9704; // @[Mux.scala 31:69:@5603.4]
  assign _T_9706 = _T_7905 ? 16'h1 : _T_9705; // @[Mux.scala 31:69:@5604.4]
  assign _T_9707 = _T_9706[0]; // @[OneHot.scala 66:30:@5605.4]
  assign _T_9708 = _T_9706[1]; // @[OneHot.scala 66:30:@5606.4]
  assign _T_9709 = _T_9706[2]; // @[OneHot.scala 66:30:@5607.4]
  assign _T_9710 = _T_9706[3]; // @[OneHot.scala 66:30:@5608.4]
  assign _T_9711 = _T_9706[4]; // @[OneHot.scala 66:30:@5609.4]
  assign _T_9712 = _T_9706[5]; // @[OneHot.scala 66:30:@5610.4]
  assign _T_9713 = _T_9706[6]; // @[OneHot.scala 66:30:@5611.4]
  assign _T_9714 = _T_9706[7]; // @[OneHot.scala 66:30:@5612.4]
  assign _T_9715 = _T_9706[8]; // @[OneHot.scala 66:30:@5613.4]
  assign _T_9716 = _T_9706[9]; // @[OneHot.scala 66:30:@5614.4]
  assign _T_9717 = _T_9706[10]; // @[OneHot.scala 66:30:@5615.4]
  assign _T_9718 = _T_9706[11]; // @[OneHot.scala 66:30:@5616.4]
  assign _T_9719 = _T_9706[12]; // @[OneHot.scala 66:30:@5617.4]
  assign _T_9720 = _T_9706[13]; // @[OneHot.scala 66:30:@5618.4]
  assign _T_9721 = _T_9706[14]; // @[OneHot.scala 66:30:@5619.4]
  assign _T_9722 = _T_9706[15]; // @[OneHot.scala 66:30:@5620.4]
  assign _T_9763 = _T_7905 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5638.4]
  assign _T_9764 = _T_7950 ? 16'h4000 : _T_9763; // @[Mux.scala 31:69:@5639.4]
  assign _T_9765 = _T_7947 ? 16'h2000 : _T_9764; // @[Mux.scala 31:69:@5640.4]
  assign _T_9766 = _T_7944 ? 16'h1000 : _T_9765; // @[Mux.scala 31:69:@5641.4]
  assign _T_9767 = _T_7941 ? 16'h800 : _T_9766; // @[Mux.scala 31:69:@5642.4]
  assign _T_9768 = _T_7938 ? 16'h400 : _T_9767; // @[Mux.scala 31:69:@5643.4]
  assign _T_9769 = _T_7935 ? 16'h200 : _T_9768; // @[Mux.scala 31:69:@5644.4]
  assign _T_9770 = _T_7932 ? 16'h100 : _T_9769; // @[Mux.scala 31:69:@5645.4]
  assign _T_9771 = _T_7929 ? 16'h80 : _T_9770; // @[Mux.scala 31:69:@5646.4]
  assign _T_9772 = _T_7926 ? 16'h40 : _T_9771; // @[Mux.scala 31:69:@5647.4]
  assign _T_9773 = _T_7923 ? 16'h20 : _T_9772; // @[Mux.scala 31:69:@5648.4]
  assign _T_9774 = _T_7920 ? 16'h10 : _T_9773; // @[Mux.scala 31:69:@5649.4]
  assign _T_9775 = _T_7917 ? 16'h8 : _T_9774; // @[Mux.scala 31:69:@5650.4]
  assign _T_9776 = _T_7914 ? 16'h4 : _T_9775; // @[Mux.scala 31:69:@5651.4]
  assign _T_9777 = _T_7911 ? 16'h2 : _T_9776; // @[Mux.scala 31:69:@5652.4]
  assign _T_9778 = _T_7908 ? 16'h1 : _T_9777; // @[Mux.scala 31:69:@5653.4]
  assign _T_9779 = _T_9778[0]; // @[OneHot.scala 66:30:@5654.4]
  assign _T_9780 = _T_9778[1]; // @[OneHot.scala 66:30:@5655.4]
  assign _T_9781 = _T_9778[2]; // @[OneHot.scala 66:30:@5656.4]
  assign _T_9782 = _T_9778[3]; // @[OneHot.scala 66:30:@5657.4]
  assign _T_9783 = _T_9778[4]; // @[OneHot.scala 66:30:@5658.4]
  assign _T_9784 = _T_9778[5]; // @[OneHot.scala 66:30:@5659.4]
  assign _T_9785 = _T_9778[6]; // @[OneHot.scala 66:30:@5660.4]
  assign _T_9786 = _T_9778[7]; // @[OneHot.scala 66:30:@5661.4]
  assign _T_9787 = _T_9778[8]; // @[OneHot.scala 66:30:@5662.4]
  assign _T_9788 = _T_9778[9]; // @[OneHot.scala 66:30:@5663.4]
  assign _T_9789 = _T_9778[10]; // @[OneHot.scala 66:30:@5664.4]
  assign _T_9790 = _T_9778[11]; // @[OneHot.scala 66:30:@5665.4]
  assign _T_9791 = _T_9778[12]; // @[OneHot.scala 66:30:@5666.4]
  assign _T_9792 = _T_9778[13]; // @[OneHot.scala 66:30:@5667.4]
  assign _T_9793 = _T_9778[14]; // @[OneHot.scala 66:30:@5668.4]
  assign _T_9794 = _T_9778[15]; // @[OneHot.scala 66:30:@5669.4]
  assign _T_9835 = _T_7908 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5687.4]
  assign _T_9836 = _T_7905 ? 16'h4000 : _T_9835; // @[Mux.scala 31:69:@5688.4]
  assign _T_9837 = _T_7950 ? 16'h2000 : _T_9836; // @[Mux.scala 31:69:@5689.4]
  assign _T_9838 = _T_7947 ? 16'h1000 : _T_9837; // @[Mux.scala 31:69:@5690.4]
  assign _T_9839 = _T_7944 ? 16'h800 : _T_9838; // @[Mux.scala 31:69:@5691.4]
  assign _T_9840 = _T_7941 ? 16'h400 : _T_9839; // @[Mux.scala 31:69:@5692.4]
  assign _T_9841 = _T_7938 ? 16'h200 : _T_9840; // @[Mux.scala 31:69:@5693.4]
  assign _T_9842 = _T_7935 ? 16'h100 : _T_9841; // @[Mux.scala 31:69:@5694.4]
  assign _T_9843 = _T_7932 ? 16'h80 : _T_9842; // @[Mux.scala 31:69:@5695.4]
  assign _T_9844 = _T_7929 ? 16'h40 : _T_9843; // @[Mux.scala 31:69:@5696.4]
  assign _T_9845 = _T_7926 ? 16'h20 : _T_9844; // @[Mux.scala 31:69:@5697.4]
  assign _T_9846 = _T_7923 ? 16'h10 : _T_9845; // @[Mux.scala 31:69:@5698.4]
  assign _T_9847 = _T_7920 ? 16'h8 : _T_9846; // @[Mux.scala 31:69:@5699.4]
  assign _T_9848 = _T_7917 ? 16'h4 : _T_9847; // @[Mux.scala 31:69:@5700.4]
  assign _T_9849 = _T_7914 ? 16'h2 : _T_9848; // @[Mux.scala 31:69:@5701.4]
  assign _T_9850 = _T_7911 ? 16'h1 : _T_9849; // @[Mux.scala 31:69:@5702.4]
  assign _T_9851 = _T_9850[0]; // @[OneHot.scala 66:30:@5703.4]
  assign _T_9852 = _T_9850[1]; // @[OneHot.scala 66:30:@5704.4]
  assign _T_9853 = _T_9850[2]; // @[OneHot.scala 66:30:@5705.4]
  assign _T_9854 = _T_9850[3]; // @[OneHot.scala 66:30:@5706.4]
  assign _T_9855 = _T_9850[4]; // @[OneHot.scala 66:30:@5707.4]
  assign _T_9856 = _T_9850[5]; // @[OneHot.scala 66:30:@5708.4]
  assign _T_9857 = _T_9850[6]; // @[OneHot.scala 66:30:@5709.4]
  assign _T_9858 = _T_9850[7]; // @[OneHot.scala 66:30:@5710.4]
  assign _T_9859 = _T_9850[8]; // @[OneHot.scala 66:30:@5711.4]
  assign _T_9860 = _T_9850[9]; // @[OneHot.scala 66:30:@5712.4]
  assign _T_9861 = _T_9850[10]; // @[OneHot.scala 66:30:@5713.4]
  assign _T_9862 = _T_9850[11]; // @[OneHot.scala 66:30:@5714.4]
  assign _T_9863 = _T_9850[12]; // @[OneHot.scala 66:30:@5715.4]
  assign _T_9864 = _T_9850[13]; // @[OneHot.scala 66:30:@5716.4]
  assign _T_9865 = _T_9850[14]; // @[OneHot.scala 66:30:@5717.4]
  assign _T_9866 = _T_9850[15]; // @[OneHot.scala 66:30:@5718.4]
  assign _T_9907 = _T_7911 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5736.4]
  assign _T_9908 = _T_7908 ? 16'h4000 : _T_9907; // @[Mux.scala 31:69:@5737.4]
  assign _T_9909 = _T_7905 ? 16'h2000 : _T_9908; // @[Mux.scala 31:69:@5738.4]
  assign _T_9910 = _T_7950 ? 16'h1000 : _T_9909; // @[Mux.scala 31:69:@5739.4]
  assign _T_9911 = _T_7947 ? 16'h800 : _T_9910; // @[Mux.scala 31:69:@5740.4]
  assign _T_9912 = _T_7944 ? 16'h400 : _T_9911; // @[Mux.scala 31:69:@5741.4]
  assign _T_9913 = _T_7941 ? 16'h200 : _T_9912; // @[Mux.scala 31:69:@5742.4]
  assign _T_9914 = _T_7938 ? 16'h100 : _T_9913; // @[Mux.scala 31:69:@5743.4]
  assign _T_9915 = _T_7935 ? 16'h80 : _T_9914; // @[Mux.scala 31:69:@5744.4]
  assign _T_9916 = _T_7932 ? 16'h40 : _T_9915; // @[Mux.scala 31:69:@5745.4]
  assign _T_9917 = _T_7929 ? 16'h20 : _T_9916; // @[Mux.scala 31:69:@5746.4]
  assign _T_9918 = _T_7926 ? 16'h10 : _T_9917; // @[Mux.scala 31:69:@5747.4]
  assign _T_9919 = _T_7923 ? 16'h8 : _T_9918; // @[Mux.scala 31:69:@5748.4]
  assign _T_9920 = _T_7920 ? 16'h4 : _T_9919; // @[Mux.scala 31:69:@5749.4]
  assign _T_9921 = _T_7917 ? 16'h2 : _T_9920; // @[Mux.scala 31:69:@5750.4]
  assign _T_9922 = _T_7914 ? 16'h1 : _T_9921; // @[Mux.scala 31:69:@5751.4]
  assign _T_9923 = _T_9922[0]; // @[OneHot.scala 66:30:@5752.4]
  assign _T_9924 = _T_9922[1]; // @[OneHot.scala 66:30:@5753.4]
  assign _T_9925 = _T_9922[2]; // @[OneHot.scala 66:30:@5754.4]
  assign _T_9926 = _T_9922[3]; // @[OneHot.scala 66:30:@5755.4]
  assign _T_9927 = _T_9922[4]; // @[OneHot.scala 66:30:@5756.4]
  assign _T_9928 = _T_9922[5]; // @[OneHot.scala 66:30:@5757.4]
  assign _T_9929 = _T_9922[6]; // @[OneHot.scala 66:30:@5758.4]
  assign _T_9930 = _T_9922[7]; // @[OneHot.scala 66:30:@5759.4]
  assign _T_9931 = _T_9922[8]; // @[OneHot.scala 66:30:@5760.4]
  assign _T_9932 = _T_9922[9]; // @[OneHot.scala 66:30:@5761.4]
  assign _T_9933 = _T_9922[10]; // @[OneHot.scala 66:30:@5762.4]
  assign _T_9934 = _T_9922[11]; // @[OneHot.scala 66:30:@5763.4]
  assign _T_9935 = _T_9922[12]; // @[OneHot.scala 66:30:@5764.4]
  assign _T_9936 = _T_9922[13]; // @[OneHot.scala 66:30:@5765.4]
  assign _T_9937 = _T_9922[14]; // @[OneHot.scala 66:30:@5766.4]
  assign _T_9938 = _T_9922[15]; // @[OneHot.scala 66:30:@5767.4]
  assign _T_9979 = _T_7914 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5785.4]
  assign _T_9980 = _T_7911 ? 16'h4000 : _T_9979; // @[Mux.scala 31:69:@5786.4]
  assign _T_9981 = _T_7908 ? 16'h2000 : _T_9980; // @[Mux.scala 31:69:@5787.4]
  assign _T_9982 = _T_7905 ? 16'h1000 : _T_9981; // @[Mux.scala 31:69:@5788.4]
  assign _T_9983 = _T_7950 ? 16'h800 : _T_9982; // @[Mux.scala 31:69:@5789.4]
  assign _T_9984 = _T_7947 ? 16'h400 : _T_9983; // @[Mux.scala 31:69:@5790.4]
  assign _T_9985 = _T_7944 ? 16'h200 : _T_9984; // @[Mux.scala 31:69:@5791.4]
  assign _T_9986 = _T_7941 ? 16'h100 : _T_9985; // @[Mux.scala 31:69:@5792.4]
  assign _T_9987 = _T_7938 ? 16'h80 : _T_9986; // @[Mux.scala 31:69:@5793.4]
  assign _T_9988 = _T_7935 ? 16'h40 : _T_9987; // @[Mux.scala 31:69:@5794.4]
  assign _T_9989 = _T_7932 ? 16'h20 : _T_9988; // @[Mux.scala 31:69:@5795.4]
  assign _T_9990 = _T_7929 ? 16'h10 : _T_9989; // @[Mux.scala 31:69:@5796.4]
  assign _T_9991 = _T_7926 ? 16'h8 : _T_9990; // @[Mux.scala 31:69:@5797.4]
  assign _T_9992 = _T_7923 ? 16'h4 : _T_9991; // @[Mux.scala 31:69:@5798.4]
  assign _T_9993 = _T_7920 ? 16'h2 : _T_9992; // @[Mux.scala 31:69:@5799.4]
  assign _T_9994 = _T_7917 ? 16'h1 : _T_9993; // @[Mux.scala 31:69:@5800.4]
  assign _T_9995 = _T_9994[0]; // @[OneHot.scala 66:30:@5801.4]
  assign _T_9996 = _T_9994[1]; // @[OneHot.scala 66:30:@5802.4]
  assign _T_9997 = _T_9994[2]; // @[OneHot.scala 66:30:@5803.4]
  assign _T_9998 = _T_9994[3]; // @[OneHot.scala 66:30:@5804.4]
  assign _T_9999 = _T_9994[4]; // @[OneHot.scala 66:30:@5805.4]
  assign _T_10000 = _T_9994[5]; // @[OneHot.scala 66:30:@5806.4]
  assign _T_10001 = _T_9994[6]; // @[OneHot.scala 66:30:@5807.4]
  assign _T_10002 = _T_9994[7]; // @[OneHot.scala 66:30:@5808.4]
  assign _T_10003 = _T_9994[8]; // @[OneHot.scala 66:30:@5809.4]
  assign _T_10004 = _T_9994[9]; // @[OneHot.scala 66:30:@5810.4]
  assign _T_10005 = _T_9994[10]; // @[OneHot.scala 66:30:@5811.4]
  assign _T_10006 = _T_9994[11]; // @[OneHot.scala 66:30:@5812.4]
  assign _T_10007 = _T_9994[12]; // @[OneHot.scala 66:30:@5813.4]
  assign _T_10008 = _T_9994[13]; // @[OneHot.scala 66:30:@5814.4]
  assign _T_10009 = _T_9994[14]; // @[OneHot.scala 66:30:@5815.4]
  assign _T_10010 = _T_9994[15]; // @[OneHot.scala 66:30:@5816.4]
  assign _T_10051 = _T_7917 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5834.4]
  assign _T_10052 = _T_7914 ? 16'h4000 : _T_10051; // @[Mux.scala 31:69:@5835.4]
  assign _T_10053 = _T_7911 ? 16'h2000 : _T_10052; // @[Mux.scala 31:69:@5836.4]
  assign _T_10054 = _T_7908 ? 16'h1000 : _T_10053; // @[Mux.scala 31:69:@5837.4]
  assign _T_10055 = _T_7905 ? 16'h800 : _T_10054; // @[Mux.scala 31:69:@5838.4]
  assign _T_10056 = _T_7950 ? 16'h400 : _T_10055; // @[Mux.scala 31:69:@5839.4]
  assign _T_10057 = _T_7947 ? 16'h200 : _T_10056; // @[Mux.scala 31:69:@5840.4]
  assign _T_10058 = _T_7944 ? 16'h100 : _T_10057; // @[Mux.scala 31:69:@5841.4]
  assign _T_10059 = _T_7941 ? 16'h80 : _T_10058; // @[Mux.scala 31:69:@5842.4]
  assign _T_10060 = _T_7938 ? 16'h40 : _T_10059; // @[Mux.scala 31:69:@5843.4]
  assign _T_10061 = _T_7935 ? 16'h20 : _T_10060; // @[Mux.scala 31:69:@5844.4]
  assign _T_10062 = _T_7932 ? 16'h10 : _T_10061; // @[Mux.scala 31:69:@5845.4]
  assign _T_10063 = _T_7929 ? 16'h8 : _T_10062; // @[Mux.scala 31:69:@5846.4]
  assign _T_10064 = _T_7926 ? 16'h4 : _T_10063; // @[Mux.scala 31:69:@5847.4]
  assign _T_10065 = _T_7923 ? 16'h2 : _T_10064; // @[Mux.scala 31:69:@5848.4]
  assign _T_10066 = _T_7920 ? 16'h1 : _T_10065; // @[Mux.scala 31:69:@5849.4]
  assign _T_10067 = _T_10066[0]; // @[OneHot.scala 66:30:@5850.4]
  assign _T_10068 = _T_10066[1]; // @[OneHot.scala 66:30:@5851.4]
  assign _T_10069 = _T_10066[2]; // @[OneHot.scala 66:30:@5852.4]
  assign _T_10070 = _T_10066[3]; // @[OneHot.scala 66:30:@5853.4]
  assign _T_10071 = _T_10066[4]; // @[OneHot.scala 66:30:@5854.4]
  assign _T_10072 = _T_10066[5]; // @[OneHot.scala 66:30:@5855.4]
  assign _T_10073 = _T_10066[6]; // @[OneHot.scala 66:30:@5856.4]
  assign _T_10074 = _T_10066[7]; // @[OneHot.scala 66:30:@5857.4]
  assign _T_10075 = _T_10066[8]; // @[OneHot.scala 66:30:@5858.4]
  assign _T_10076 = _T_10066[9]; // @[OneHot.scala 66:30:@5859.4]
  assign _T_10077 = _T_10066[10]; // @[OneHot.scala 66:30:@5860.4]
  assign _T_10078 = _T_10066[11]; // @[OneHot.scala 66:30:@5861.4]
  assign _T_10079 = _T_10066[12]; // @[OneHot.scala 66:30:@5862.4]
  assign _T_10080 = _T_10066[13]; // @[OneHot.scala 66:30:@5863.4]
  assign _T_10081 = _T_10066[14]; // @[OneHot.scala 66:30:@5864.4]
  assign _T_10082 = _T_10066[15]; // @[OneHot.scala 66:30:@5865.4]
  assign _T_10123 = _T_7920 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5883.4]
  assign _T_10124 = _T_7917 ? 16'h4000 : _T_10123; // @[Mux.scala 31:69:@5884.4]
  assign _T_10125 = _T_7914 ? 16'h2000 : _T_10124; // @[Mux.scala 31:69:@5885.4]
  assign _T_10126 = _T_7911 ? 16'h1000 : _T_10125; // @[Mux.scala 31:69:@5886.4]
  assign _T_10127 = _T_7908 ? 16'h800 : _T_10126; // @[Mux.scala 31:69:@5887.4]
  assign _T_10128 = _T_7905 ? 16'h400 : _T_10127; // @[Mux.scala 31:69:@5888.4]
  assign _T_10129 = _T_7950 ? 16'h200 : _T_10128; // @[Mux.scala 31:69:@5889.4]
  assign _T_10130 = _T_7947 ? 16'h100 : _T_10129; // @[Mux.scala 31:69:@5890.4]
  assign _T_10131 = _T_7944 ? 16'h80 : _T_10130; // @[Mux.scala 31:69:@5891.4]
  assign _T_10132 = _T_7941 ? 16'h40 : _T_10131; // @[Mux.scala 31:69:@5892.4]
  assign _T_10133 = _T_7938 ? 16'h20 : _T_10132; // @[Mux.scala 31:69:@5893.4]
  assign _T_10134 = _T_7935 ? 16'h10 : _T_10133; // @[Mux.scala 31:69:@5894.4]
  assign _T_10135 = _T_7932 ? 16'h8 : _T_10134; // @[Mux.scala 31:69:@5895.4]
  assign _T_10136 = _T_7929 ? 16'h4 : _T_10135; // @[Mux.scala 31:69:@5896.4]
  assign _T_10137 = _T_7926 ? 16'h2 : _T_10136; // @[Mux.scala 31:69:@5897.4]
  assign _T_10138 = _T_7923 ? 16'h1 : _T_10137; // @[Mux.scala 31:69:@5898.4]
  assign _T_10139 = _T_10138[0]; // @[OneHot.scala 66:30:@5899.4]
  assign _T_10140 = _T_10138[1]; // @[OneHot.scala 66:30:@5900.4]
  assign _T_10141 = _T_10138[2]; // @[OneHot.scala 66:30:@5901.4]
  assign _T_10142 = _T_10138[3]; // @[OneHot.scala 66:30:@5902.4]
  assign _T_10143 = _T_10138[4]; // @[OneHot.scala 66:30:@5903.4]
  assign _T_10144 = _T_10138[5]; // @[OneHot.scala 66:30:@5904.4]
  assign _T_10145 = _T_10138[6]; // @[OneHot.scala 66:30:@5905.4]
  assign _T_10146 = _T_10138[7]; // @[OneHot.scala 66:30:@5906.4]
  assign _T_10147 = _T_10138[8]; // @[OneHot.scala 66:30:@5907.4]
  assign _T_10148 = _T_10138[9]; // @[OneHot.scala 66:30:@5908.4]
  assign _T_10149 = _T_10138[10]; // @[OneHot.scala 66:30:@5909.4]
  assign _T_10150 = _T_10138[11]; // @[OneHot.scala 66:30:@5910.4]
  assign _T_10151 = _T_10138[12]; // @[OneHot.scala 66:30:@5911.4]
  assign _T_10152 = _T_10138[13]; // @[OneHot.scala 66:30:@5912.4]
  assign _T_10153 = _T_10138[14]; // @[OneHot.scala 66:30:@5913.4]
  assign _T_10154 = _T_10138[15]; // @[OneHot.scala 66:30:@5914.4]
  assign _T_10195 = _T_7923 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5932.4]
  assign _T_10196 = _T_7920 ? 16'h4000 : _T_10195; // @[Mux.scala 31:69:@5933.4]
  assign _T_10197 = _T_7917 ? 16'h2000 : _T_10196; // @[Mux.scala 31:69:@5934.4]
  assign _T_10198 = _T_7914 ? 16'h1000 : _T_10197; // @[Mux.scala 31:69:@5935.4]
  assign _T_10199 = _T_7911 ? 16'h800 : _T_10198; // @[Mux.scala 31:69:@5936.4]
  assign _T_10200 = _T_7908 ? 16'h400 : _T_10199; // @[Mux.scala 31:69:@5937.4]
  assign _T_10201 = _T_7905 ? 16'h200 : _T_10200; // @[Mux.scala 31:69:@5938.4]
  assign _T_10202 = _T_7950 ? 16'h100 : _T_10201; // @[Mux.scala 31:69:@5939.4]
  assign _T_10203 = _T_7947 ? 16'h80 : _T_10202; // @[Mux.scala 31:69:@5940.4]
  assign _T_10204 = _T_7944 ? 16'h40 : _T_10203; // @[Mux.scala 31:69:@5941.4]
  assign _T_10205 = _T_7941 ? 16'h20 : _T_10204; // @[Mux.scala 31:69:@5942.4]
  assign _T_10206 = _T_7938 ? 16'h10 : _T_10205; // @[Mux.scala 31:69:@5943.4]
  assign _T_10207 = _T_7935 ? 16'h8 : _T_10206; // @[Mux.scala 31:69:@5944.4]
  assign _T_10208 = _T_7932 ? 16'h4 : _T_10207; // @[Mux.scala 31:69:@5945.4]
  assign _T_10209 = _T_7929 ? 16'h2 : _T_10208; // @[Mux.scala 31:69:@5946.4]
  assign _T_10210 = _T_7926 ? 16'h1 : _T_10209; // @[Mux.scala 31:69:@5947.4]
  assign _T_10211 = _T_10210[0]; // @[OneHot.scala 66:30:@5948.4]
  assign _T_10212 = _T_10210[1]; // @[OneHot.scala 66:30:@5949.4]
  assign _T_10213 = _T_10210[2]; // @[OneHot.scala 66:30:@5950.4]
  assign _T_10214 = _T_10210[3]; // @[OneHot.scala 66:30:@5951.4]
  assign _T_10215 = _T_10210[4]; // @[OneHot.scala 66:30:@5952.4]
  assign _T_10216 = _T_10210[5]; // @[OneHot.scala 66:30:@5953.4]
  assign _T_10217 = _T_10210[6]; // @[OneHot.scala 66:30:@5954.4]
  assign _T_10218 = _T_10210[7]; // @[OneHot.scala 66:30:@5955.4]
  assign _T_10219 = _T_10210[8]; // @[OneHot.scala 66:30:@5956.4]
  assign _T_10220 = _T_10210[9]; // @[OneHot.scala 66:30:@5957.4]
  assign _T_10221 = _T_10210[10]; // @[OneHot.scala 66:30:@5958.4]
  assign _T_10222 = _T_10210[11]; // @[OneHot.scala 66:30:@5959.4]
  assign _T_10223 = _T_10210[12]; // @[OneHot.scala 66:30:@5960.4]
  assign _T_10224 = _T_10210[13]; // @[OneHot.scala 66:30:@5961.4]
  assign _T_10225 = _T_10210[14]; // @[OneHot.scala 66:30:@5962.4]
  assign _T_10226 = _T_10210[15]; // @[OneHot.scala 66:30:@5963.4]
  assign _T_10267 = _T_7926 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@5981.4]
  assign _T_10268 = _T_7923 ? 16'h4000 : _T_10267; // @[Mux.scala 31:69:@5982.4]
  assign _T_10269 = _T_7920 ? 16'h2000 : _T_10268; // @[Mux.scala 31:69:@5983.4]
  assign _T_10270 = _T_7917 ? 16'h1000 : _T_10269; // @[Mux.scala 31:69:@5984.4]
  assign _T_10271 = _T_7914 ? 16'h800 : _T_10270; // @[Mux.scala 31:69:@5985.4]
  assign _T_10272 = _T_7911 ? 16'h400 : _T_10271; // @[Mux.scala 31:69:@5986.4]
  assign _T_10273 = _T_7908 ? 16'h200 : _T_10272; // @[Mux.scala 31:69:@5987.4]
  assign _T_10274 = _T_7905 ? 16'h100 : _T_10273; // @[Mux.scala 31:69:@5988.4]
  assign _T_10275 = _T_7950 ? 16'h80 : _T_10274; // @[Mux.scala 31:69:@5989.4]
  assign _T_10276 = _T_7947 ? 16'h40 : _T_10275; // @[Mux.scala 31:69:@5990.4]
  assign _T_10277 = _T_7944 ? 16'h20 : _T_10276; // @[Mux.scala 31:69:@5991.4]
  assign _T_10278 = _T_7941 ? 16'h10 : _T_10277; // @[Mux.scala 31:69:@5992.4]
  assign _T_10279 = _T_7938 ? 16'h8 : _T_10278; // @[Mux.scala 31:69:@5993.4]
  assign _T_10280 = _T_7935 ? 16'h4 : _T_10279; // @[Mux.scala 31:69:@5994.4]
  assign _T_10281 = _T_7932 ? 16'h2 : _T_10280; // @[Mux.scala 31:69:@5995.4]
  assign _T_10282 = _T_7929 ? 16'h1 : _T_10281; // @[Mux.scala 31:69:@5996.4]
  assign _T_10283 = _T_10282[0]; // @[OneHot.scala 66:30:@5997.4]
  assign _T_10284 = _T_10282[1]; // @[OneHot.scala 66:30:@5998.4]
  assign _T_10285 = _T_10282[2]; // @[OneHot.scala 66:30:@5999.4]
  assign _T_10286 = _T_10282[3]; // @[OneHot.scala 66:30:@6000.4]
  assign _T_10287 = _T_10282[4]; // @[OneHot.scala 66:30:@6001.4]
  assign _T_10288 = _T_10282[5]; // @[OneHot.scala 66:30:@6002.4]
  assign _T_10289 = _T_10282[6]; // @[OneHot.scala 66:30:@6003.4]
  assign _T_10290 = _T_10282[7]; // @[OneHot.scala 66:30:@6004.4]
  assign _T_10291 = _T_10282[8]; // @[OneHot.scala 66:30:@6005.4]
  assign _T_10292 = _T_10282[9]; // @[OneHot.scala 66:30:@6006.4]
  assign _T_10293 = _T_10282[10]; // @[OneHot.scala 66:30:@6007.4]
  assign _T_10294 = _T_10282[11]; // @[OneHot.scala 66:30:@6008.4]
  assign _T_10295 = _T_10282[12]; // @[OneHot.scala 66:30:@6009.4]
  assign _T_10296 = _T_10282[13]; // @[OneHot.scala 66:30:@6010.4]
  assign _T_10297 = _T_10282[14]; // @[OneHot.scala 66:30:@6011.4]
  assign _T_10298 = _T_10282[15]; // @[OneHot.scala 66:30:@6012.4]
  assign _T_10339 = _T_7929 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6030.4]
  assign _T_10340 = _T_7926 ? 16'h4000 : _T_10339; // @[Mux.scala 31:69:@6031.4]
  assign _T_10341 = _T_7923 ? 16'h2000 : _T_10340; // @[Mux.scala 31:69:@6032.4]
  assign _T_10342 = _T_7920 ? 16'h1000 : _T_10341; // @[Mux.scala 31:69:@6033.4]
  assign _T_10343 = _T_7917 ? 16'h800 : _T_10342; // @[Mux.scala 31:69:@6034.4]
  assign _T_10344 = _T_7914 ? 16'h400 : _T_10343; // @[Mux.scala 31:69:@6035.4]
  assign _T_10345 = _T_7911 ? 16'h200 : _T_10344; // @[Mux.scala 31:69:@6036.4]
  assign _T_10346 = _T_7908 ? 16'h100 : _T_10345; // @[Mux.scala 31:69:@6037.4]
  assign _T_10347 = _T_7905 ? 16'h80 : _T_10346; // @[Mux.scala 31:69:@6038.4]
  assign _T_10348 = _T_7950 ? 16'h40 : _T_10347; // @[Mux.scala 31:69:@6039.4]
  assign _T_10349 = _T_7947 ? 16'h20 : _T_10348; // @[Mux.scala 31:69:@6040.4]
  assign _T_10350 = _T_7944 ? 16'h10 : _T_10349; // @[Mux.scala 31:69:@6041.4]
  assign _T_10351 = _T_7941 ? 16'h8 : _T_10350; // @[Mux.scala 31:69:@6042.4]
  assign _T_10352 = _T_7938 ? 16'h4 : _T_10351; // @[Mux.scala 31:69:@6043.4]
  assign _T_10353 = _T_7935 ? 16'h2 : _T_10352; // @[Mux.scala 31:69:@6044.4]
  assign _T_10354 = _T_7932 ? 16'h1 : _T_10353; // @[Mux.scala 31:69:@6045.4]
  assign _T_10355 = _T_10354[0]; // @[OneHot.scala 66:30:@6046.4]
  assign _T_10356 = _T_10354[1]; // @[OneHot.scala 66:30:@6047.4]
  assign _T_10357 = _T_10354[2]; // @[OneHot.scala 66:30:@6048.4]
  assign _T_10358 = _T_10354[3]; // @[OneHot.scala 66:30:@6049.4]
  assign _T_10359 = _T_10354[4]; // @[OneHot.scala 66:30:@6050.4]
  assign _T_10360 = _T_10354[5]; // @[OneHot.scala 66:30:@6051.4]
  assign _T_10361 = _T_10354[6]; // @[OneHot.scala 66:30:@6052.4]
  assign _T_10362 = _T_10354[7]; // @[OneHot.scala 66:30:@6053.4]
  assign _T_10363 = _T_10354[8]; // @[OneHot.scala 66:30:@6054.4]
  assign _T_10364 = _T_10354[9]; // @[OneHot.scala 66:30:@6055.4]
  assign _T_10365 = _T_10354[10]; // @[OneHot.scala 66:30:@6056.4]
  assign _T_10366 = _T_10354[11]; // @[OneHot.scala 66:30:@6057.4]
  assign _T_10367 = _T_10354[12]; // @[OneHot.scala 66:30:@6058.4]
  assign _T_10368 = _T_10354[13]; // @[OneHot.scala 66:30:@6059.4]
  assign _T_10369 = _T_10354[14]; // @[OneHot.scala 66:30:@6060.4]
  assign _T_10370 = _T_10354[15]; // @[OneHot.scala 66:30:@6061.4]
  assign _T_10411 = _T_7932 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6079.4]
  assign _T_10412 = _T_7929 ? 16'h4000 : _T_10411; // @[Mux.scala 31:69:@6080.4]
  assign _T_10413 = _T_7926 ? 16'h2000 : _T_10412; // @[Mux.scala 31:69:@6081.4]
  assign _T_10414 = _T_7923 ? 16'h1000 : _T_10413; // @[Mux.scala 31:69:@6082.4]
  assign _T_10415 = _T_7920 ? 16'h800 : _T_10414; // @[Mux.scala 31:69:@6083.4]
  assign _T_10416 = _T_7917 ? 16'h400 : _T_10415; // @[Mux.scala 31:69:@6084.4]
  assign _T_10417 = _T_7914 ? 16'h200 : _T_10416; // @[Mux.scala 31:69:@6085.4]
  assign _T_10418 = _T_7911 ? 16'h100 : _T_10417; // @[Mux.scala 31:69:@6086.4]
  assign _T_10419 = _T_7908 ? 16'h80 : _T_10418; // @[Mux.scala 31:69:@6087.4]
  assign _T_10420 = _T_7905 ? 16'h40 : _T_10419; // @[Mux.scala 31:69:@6088.4]
  assign _T_10421 = _T_7950 ? 16'h20 : _T_10420; // @[Mux.scala 31:69:@6089.4]
  assign _T_10422 = _T_7947 ? 16'h10 : _T_10421; // @[Mux.scala 31:69:@6090.4]
  assign _T_10423 = _T_7944 ? 16'h8 : _T_10422; // @[Mux.scala 31:69:@6091.4]
  assign _T_10424 = _T_7941 ? 16'h4 : _T_10423; // @[Mux.scala 31:69:@6092.4]
  assign _T_10425 = _T_7938 ? 16'h2 : _T_10424; // @[Mux.scala 31:69:@6093.4]
  assign _T_10426 = _T_7935 ? 16'h1 : _T_10425; // @[Mux.scala 31:69:@6094.4]
  assign _T_10427 = _T_10426[0]; // @[OneHot.scala 66:30:@6095.4]
  assign _T_10428 = _T_10426[1]; // @[OneHot.scala 66:30:@6096.4]
  assign _T_10429 = _T_10426[2]; // @[OneHot.scala 66:30:@6097.4]
  assign _T_10430 = _T_10426[3]; // @[OneHot.scala 66:30:@6098.4]
  assign _T_10431 = _T_10426[4]; // @[OneHot.scala 66:30:@6099.4]
  assign _T_10432 = _T_10426[5]; // @[OneHot.scala 66:30:@6100.4]
  assign _T_10433 = _T_10426[6]; // @[OneHot.scala 66:30:@6101.4]
  assign _T_10434 = _T_10426[7]; // @[OneHot.scala 66:30:@6102.4]
  assign _T_10435 = _T_10426[8]; // @[OneHot.scala 66:30:@6103.4]
  assign _T_10436 = _T_10426[9]; // @[OneHot.scala 66:30:@6104.4]
  assign _T_10437 = _T_10426[10]; // @[OneHot.scala 66:30:@6105.4]
  assign _T_10438 = _T_10426[11]; // @[OneHot.scala 66:30:@6106.4]
  assign _T_10439 = _T_10426[12]; // @[OneHot.scala 66:30:@6107.4]
  assign _T_10440 = _T_10426[13]; // @[OneHot.scala 66:30:@6108.4]
  assign _T_10441 = _T_10426[14]; // @[OneHot.scala 66:30:@6109.4]
  assign _T_10442 = _T_10426[15]; // @[OneHot.scala 66:30:@6110.4]
  assign _T_10483 = _T_7935 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6128.4]
  assign _T_10484 = _T_7932 ? 16'h4000 : _T_10483; // @[Mux.scala 31:69:@6129.4]
  assign _T_10485 = _T_7929 ? 16'h2000 : _T_10484; // @[Mux.scala 31:69:@6130.4]
  assign _T_10486 = _T_7926 ? 16'h1000 : _T_10485; // @[Mux.scala 31:69:@6131.4]
  assign _T_10487 = _T_7923 ? 16'h800 : _T_10486; // @[Mux.scala 31:69:@6132.4]
  assign _T_10488 = _T_7920 ? 16'h400 : _T_10487; // @[Mux.scala 31:69:@6133.4]
  assign _T_10489 = _T_7917 ? 16'h200 : _T_10488; // @[Mux.scala 31:69:@6134.4]
  assign _T_10490 = _T_7914 ? 16'h100 : _T_10489; // @[Mux.scala 31:69:@6135.4]
  assign _T_10491 = _T_7911 ? 16'h80 : _T_10490; // @[Mux.scala 31:69:@6136.4]
  assign _T_10492 = _T_7908 ? 16'h40 : _T_10491; // @[Mux.scala 31:69:@6137.4]
  assign _T_10493 = _T_7905 ? 16'h20 : _T_10492; // @[Mux.scala 31:69:@6138.4]
  assign _T_10494 = _T_7950 ? 16'h10 : _T_10493; // @[Mux.scala 31:69:@6139.4]
  assign _T_10495 = _T_7947 ? 16'h8 : _T_10494; // @[Mux.scala 31:69:@6140.4]
  assign _T_10496 = _T_7944 ? 16'h4 : _T_10495; // @[Mux.scala 31:69:@6141.4]
  assign _T_10497 = _T_7941 ? 16'h2 : _T_10496; // @[Mux.scala 31:69:@6142.4]
  assign _T_10498 = _T_7938 ? 16'h1 : _T_10497; // @[Mux.scala 31:69:@6143.4]
  assign _T_10499 = _T_10498[0]; // @[OneHot.scala 66:30:@6144.4]
  assign _T_10500 = _T_10498[1]; // @[OneHot.scala 66:30:@6145.4]
  assign _T_10501 = _T_10498[2]; // @[OneHot.scala 66:30:@6146.4]
  assign _T_10502 = _T_10498[3]; // @[OneHot.scala 66:30:@6147.4]
  assign _T_10503 = _T_10498[4]; // @[OneHot.scala 66:30:@6148.4]
  assign _T_10504 = _T_10498[5]; // @[OneHot.scala 66:30:@6149.4]
  assign _T_10505 = _T_10498[6]; // @[OneHot.scala 66:30:@6150.4]
  assign _T_10506 = _T_10498[7]; // @[OneHot.scala 66:30:@6151.4]
  assign _T_10507 = _T_10498[8]; // @[OneHot.scala 66:30:@6152.4]
  assign _T_10508 = _T_10498[9]; // @[OneHot.scala 66:30:@6153.4]
  assign _T_10509 = _T_10498[10]; // @[OneHot.scala 66:30:@6154.4]
  assign _T_10510 = _T_10498[11]; // @[OneHot.scala 66:30:@6155.4]
  assign _T_10511 = _T_10498[12]; // @[OneHot.scala 66:30:@6156.4]
  assign _T_10512 = _T_10498[13]; // @[OneHot.scala 66:30:@6157.4]
  assign _T_10513 = _T_10498[14]; // @[OneHot.scala 66:30:@6158.4]
  assign _T_10514 = _T_10498[15]; // @[OneHot.scala 66:30:@6159.4]
  assign _T_10555 = _T_7938 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6177.4]
  assign _T_10556 = _T_7935 ? 16'h4000 : _T_10555; // @[Mux.scala 31:69:@6178.4]
  assign _T_10557 = _T_7932 ? 16'h2000 : _T_10556; // @[Mux.scala 31:69:@6179.4]
  assign _T_10558 = _T_7929 ? 16'h1000 : _T_10557; // @[Mux.scala 31:69:@6180.4]
  assign _T_10559 = _T_7926 ? 16'h800 : _T_10558; // @[Mux.scala 31:69:@6181.4]
  assign _T_10560 = _T_7923 ? 16'h400 : _T_10559; // @[Mux.scala 31:69:@6182.4]
  assign _T_10561 = _T_7920 ? 16'h200 : _T_10560; // @[Mux.scala 31:69:@6183.4]
  assign _T_10562 = _T_7917 ? 16'h100 : _T_10561; // @[Mux.scala 31:69:@6184.4]
  assign _T_10563 = _T_7914 ? 16'h80 : _T_10562; // @[Mux.scala 31:69:@6185.4]
  assign _T_10564 = _T_7911 ? 16'h40 : _T_10563; // @[Mux.scala 31:69:@6186.4]
  assign _T_10565 = _T_7908 ? 16'h20 : _T_10564; // @[Mux.scala 31:69:@6187.4]
  assign _T_10566 = _T_7905 ? 16'h10 : _T_10565; // @[Mux.scala 31:69:@6188.4]
  assign _T_10567 = _T_7950 ? 16'h8 : _T_10566; // @[Mux.scala 31:69:@6189.4]
  assign _T_10568 = _T_7947 ? 16'h4 : _T_10567; // @[Mux.scala 31:69:@6190.4]
  assign _T_10569 = _T_7944 ? 16'h2 : _T_10568; // @[Mux.scala 31:69:@6191.4]
  assign _T_10570 = _T_7941 ? 16'h1 : _T_10569; // @[Mux.scala 31:69:@6192.4]
  assign _T_10571 = _T_10570[0]; // @[OneHot.scala 66:30:@6193.4]
  assign _T_10572 = _T_10570[1]; // @[OneHot.scala 66:30:@6194.4]
  assign _T_10573 = _T_10570[2]; // @[OneHot.scala 66:30:@6195.4]
  assign _T_10574 = _T_10570[3]; // @[OneHot.scala 66:30:@6196.4]
  assign _T_10575 = _T_10570[4]; // @[OneHot.scala 66:30:@6197.4]
  assign _T_10576 = _T_10570[5]; // @[OneHot.scala 66:30:@6198.4]
  assign _T_10577 = _T_10570[6]; // @[OneHot.scala 66:30:@6199.4]
  assign _T_10578 = _T_10570[7]; // @[OneHot.scala 66:30:@6200.4]
  assign _T_10579 = _T_10570[8]; // @[OneHot.scala 66:30:@6201.4]
  assign _T_10580 = _T_10570[9]; // @[OneHot.scala 66:30:@6202.4]
  assign _T_10581 = _T_10570[10]; // @[OneHot.scala 66:30:@6203.4]
  assign _T_10582 = _T_10570[11]; // @[OneHot.scala 66:30:@6204.4]
  assign _T_10583 = _T_10570[12]; // @[OneHot.scala 66:30:@6205.4]
  assign _T_10584 = _T_10570[13]; // @[OneHot.scala 66:30:@6206.4]
  assign _T_10585 = _T_10570[14]; // @[OneHot.scala 66:30:@6207.4]
  assign _T_10586 = _T_10570[15]; // @[OneHot.scala 66:30:@6208.4]
  assign _T_10627 = _T_7941 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6226.4]
  assign _T_10628 = _T_7938 ? 16'h4000 : _T_10627; // @[Mux.scala 31:69:@6227.4]
  assign _T_10629 = _T_7935 ? 16'h2000 : _T_10628; // @[Mux.scala 31:69:@6228.4]
  assign _T_10630 = _T_7932 ? 16'h1000 : _T_10629; // @[Mux.scala 31:69:@6229.4]
  assign _T_10631 = _T_7929 ? 16'h800 : _T_10630; // @[Mux.scala 31:69:@6230.4]
  assign _T_10632 = _T_7926 ? 16'h400 : _T_10631; // @[Mux.scala 31:69:@6231.4]
  assign _T_10633 = _T_7923 ? 16'h200 : _T_10632; // @[Mux.scala 31:69:@6232.4]
  assign _T_10634 = _T_7920 ? 16'h100 : _T_10633; // @[Mux.scala 31:69:@6233.4]
  assign _T_10635 = _T_7917 ? 16'h80 : _T_10634; // @[Mux.scala 31:69:@6234.4]
  assign _T_10636 = _T_7914 ? 16'h40 : _T_10635; // @[Mux.scala 31:69:@6235.4]
  assign _T_10637 = _T_7911 ? 16'h20 : _T_10636; // @[Mux.scala 31:69:@6236.4]
  assign _T_10638 = _T_7908 ? 16'h10 : _T_10637; // @[Mux.scala 31:69:@6237.4]
  assign _T_10639 = _T_7905 ? 16'h8 : _T_10638; // @[Mux.scala 31:69:@6238.4]
  assign _T_10640 = _T_7950 ? 16'h4 : _T_10639; // @[Mux.scala 31:69:@6239.4]
  assign _T_10641 = _T_7947 ? 16'h2 : _T_10640; // @[Mux.scala 31:69:@6240.4]
  assign _T_10642 = _T_7944 ? 16'h1 : _T_10641; // @[Mux.scala 31:69:@6241.4]
  assign _T_10643 = _T_10642[0]; // @[OneHot.scala 66:30:@6242.4]
  assign _T_10644 = _T_10642[1]; // @[OneHot.scala 66:30:@6243.4]
  assign _T_10645 = _T_10642[2]; // @[OneHot.scala 66:30:@6244.4]
  assign _T_10646 = _T_10642[3]; // @[OneHot.scala 66:30:@6245.4]
  assign _T_10647 = _T_10642[4]; // @[OneHot.scala 66:30:@6246.4]
  assign _T_10648 = _T_10642[5]; // @[OneHot.scala 66:30:@6247.4]
  assign _T_10649 = _T_10642[6]; // @[OneHot.scala 66:30:@6248.4]
  assign _T_10650 = _T_10642[7]; // @[OneHot.scala 66:30:@6249.4]
  assign _T_10651 = _T_10642[8]; // @[OneHot.scala 66:30:@6250.4]
  assign _T_10652 = _T_10642[9]; // @[OneHot.scala 66:30:@6251.4]
  assign _T_10653 = _T_10642[10]; // @[OneHot.scala 66:30:@6252.4]
  assign _T_10654 = _T_10642[11]; // @[OneHot.scala 66:30:@6253.4]
  assign _T_10655 = _T_10642[12]; // @[OneHot.scala 66:30:@6254.4]
  assign _T_10656 = _T_10642[13]; // @[OneHot.scala 66:30:@6255.4]
  assign _T_10657 = _T_10642[14]; // @[OneHot.scala 66:30:@6256.4]
  assign _T_10658 = _T_10642[15]; // @[OneHot.scala 66:30:@6257.4]
  assign _T_10699 = _T_7944 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6275.4]
  assign _T_10700 = _T_7941 ? 16'h4000 : _T_10699; // @[Mux.scala 31:69:@6276.4]
  assign _T_10701 = _T_7938 ? 16'h2000 : _T_10700; // @[Mux.scala 31:69:@6277.4]
  assign _T_10702 = _T_7935 ? 16'h1000 : _T_10701; // @[Mux.scala 31:69:@6278.4]
  assign _T_10703 = _T_7932 ? 16'h800 : _T_10702; // @[Mux.scala 31:69:@6279.4]
  assign _T_10704 = _T_7929 ? 16'h400 : _T_10703; // @[Mux.scala 31:69:@6280.4]
  assign _T_10705 = _T_7926 ? 16'h200 : _T_10704; // @[Mux.scala 31:69:@6281.4]
  assign _T_10706 = _T_7923 ? 16'h100 : _T_10705; // @[Mux.scala 31:69:@6282.4]
  assign _T_10707 = _T_7920 ? 16'h80 : _T_10706; // @[Mux.scala 31:69:@6283.4]
  assign _T_10708 = _T_7917 ? 16'h40 : _T_10707; // @[Mux.scala 31:69:@6284.4]
  assign _T_10709 = _T_7914 ? 16'h20 : _T_10708; // @[Mux.scala 31:69:@6285.4]
  assign _T_10710 = _T_7911 ? 16'h10 : _T_10709; // @[Mux.scala 31:69:@6286.4]
  assign _T_10711 = _T_7908 ? 16'h8 : _T_10710; // @[Mux.scala 31:69:@6287.4]
  assign _T_10712 = _T_7905 ? 16'h4 : _T_10711; // @[Mux.scala 31:69:@6288.4]
  assign _T_10713 = _T_7950 ? 16'h2 : _T_10712; // @[Mux.scala 31:69:@6289.4]
  assign _T_10714 = _T_7947 ? 16'h1 : _T_10713; // @[Mux.scala 31:69:@6290.4]
  assign _T_10715 = _T_10714[0]; // @[OneHot.scala 66:30:@6291.4]
  assign _T_10716 = _T_10714[1]; // @[OneHot.scala 66:30:@6292.4]
  assign _T_10717 = _T_10714[2]; // @[OneHot.scala 66:30:@6293.4]
  assign _T_10718 = _T_10714[3]; // @[OneHot.scala 66:30:@6294.4]
  assign _T_10719 = _T_10714[4]; // @[OneHot.scala 66:30:@6295.4]
  assign _T_10720 = _T_10714[5]; // @[OneHot.scala 66:30:@6296.4]
  assign _T_10721 = _T_10714[6]; // @[OneHot.scala 66:30:@6297.4]
  assign _T_10722 = _T_10714[7]; // @[OneHot.scala 66:30:@6298.4]
  assign _T_10723 = _T_10714[8]; // @[OneHot.scala 66:30:@6299.4]
  assign _T_10724 = _T_10714[9]; // @[OneHot.scala 66:30:@6300.4]
  assign _T_10725 = _T_10714[10]; // @[OneHot.scala 66:30:@6301.4]
  assign _T_10726 = _T_10714[11]; // @[OneHot.scala 66:30:@6302.4]
  assign _T_10727 = _T_10714[12]; // @[OneHot.scala 66:30:@6303.4]
  assign _T_10728 = _T_10714[13]; // @[OneHot.scala 66:30:@6304.4]
  assign _T_10729 = _T_10714[14]; // @[OneHot.scala 66:30:@6305.4]
  assign _T_10730 = _T_10714[15]; // @[OneHot.scala 66:30:@6306.4]
  assign _T_10771 = _T_7947 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@6324.4]
  assign _T_10772 = _T_7944 ? 16'h4000 : _T_10771; // @[Mux.scala 31:69:@6325.4]
  assign _T_10773 = _T_7941 ? 16'h2000 : _T_10772; // @[Mux.scala 31:69:@6326.4]
  assign _T_10774 = _T_7938 ? 16'h1000 : _T_10773; // @[Mux.scala 31:69:@6327.4]
  assign _T_10775 = _T_7935 ? 16'h800 : _T_10774; // @[Mux.scala 31:69:@6328.4]
  assign _T_10776 = _T_7932 ? 16'h400 : _T_10775; // @[Mux.scala 31:69:@6329.4]
  assign _T_10777 = _T_7929 ? 16'h200 : _T_10776; // @[Mux.scala 31:69:@6330.4]
  assign _T_10778 = _T_7926 ? 16'h100 : _T_10777; // @[Mux.scala 31:69:@6331.4]
  assign _T_10779 = _T_7923 ? 16'h80 : _T_10778; // @[Mux.scala 31:69:@6332.4]
  assign _T_10780 = _T_7920 ? 16'h40 : _T_10779; // @[Mux.scala 31:69:@6333.4]
  assign _T_10781 = _T_7917 ? 16'h20 : _T_10780; // @[Mux.scala 31:69:@6334.4]
  assign _T_10782 = _T_7914 ? 16'h10 : _T_10781; // @[Mux.scala 31:69:@6335.4]
  assign _T_10783 = _T_7911 ? 16'h8 : _T_10782; // @[Mux.scala 31:69:@6336.4]
  assign _T_10784 = _T_7908 ? 16'h4 : _T_10783; // @[Mux.scala 31:69:@6337.4]
  assign _T_10785 = _T_7905 ? 16'h2 : _T_10784; // @[Mux.scala 31:69:@6338.4]
  assign _T_10786 = _T_7950 ? 16'h1 : _T_10785; // @[Mux.scala 31:69:@6339.4]
  assign _T_10787 = _T_10786[0]; // @[OneHot.scala 66:30:@6340.4]
  assign _T_10788 = _T_10786[1]; // @[OneHot.scala 66:30:@6341.4]
  assign _T_10789 = _T_10786[2]; // @[OneHot.scala 66:30:@6342.4]
  assign _T_10790 = _T_10786[3]; // @[OneHot.scala 66:30:@6343.4]
  assign _T_10791 = _T_10786[4]; // @[OneHot.scala 66:30:@6344.4]
  assign _T_10792 = _T_10786[5]; // @[OneHot.scala 66:30:@6345.4]
  assign _T_10793 = _T_10786[6]; // @[OneHot.scala 66:30:@6346.4]
  assign _T_10794 = _T_10786[7]; // @[OneHot.scala 66:30:@6347.4]
  assign _T_10795 = _T_10786[8]; // @[OneHot.scala 66:30:@6348.4]
  assign _T_10796 = _T_10786[9]; // @[OneHot.scala 66:30:@6349.4]
  assign _T_10797 = _T_10786[10]; // @[OneHot.scala 66:30:@6350.4]
  assign _T_10798 = _T_10786[11]; // @[OneHot.scala 66:30:@6351.4]
  assign _T_10799 = _T_10786[12]; // @[OneHot.scala 66:30:@6352.4]
  assign _T_10800 = _T_10786[13]; // @[OneHot.scala 66:30:@6353.4]
  assign _T_10801 = _T_10786[14]; // @[OneHot.scala 66:30:@6354.4]
  assign _T_10802 = _T_10786[15]; // @[OneHot.scala 66:30:@6355.4]
  assign _T_10867 = {_T_9714,_T_9713,_T_9712,_T_9711,_T_9710,_T_9709,_T_9708,_T_9707}; // @[Mux.scala 19:72:@6379.4]
  assign _T_10875 = {_T_9722,_T_9721,_T_9720,_T_9719,_T_9718,_T_9717,_T_9716,_T_9715,_T_10867}; // @[Mux.scala 19:72:@6387.4]
  assign _T_10877 = _T_4521 ? _T_10875 : 16'h0; // @[Mux.scala 19:72:@6388.4]
  assign _T_10884 = {_T_9785,_T_9784,_T_9783,_T_9782,_T_9781,_T_9780,_T_9779,_T_9794}; // @[Mux.scala 19:72:@6395.4]
  assign _T_10892 = {_T_9793,_T_9792,_T_9791,_T_9790,_T_9789,_T_9788,_T_9787,_T_9786,_T_10884}; // @[Mux.scala 19:72:@6403.4]
  assign _T_10894 = _T_4522 ? _T_10892 : 16'h0; // @[Mux.scala 19:72:@6404.4]
  assign _T_10901 = {_T_9856,_T_9855,_T_9854,_T_9853,_T_9852,_T_9851,_T_9866,_T_9865}; // @[Mux.scala 19:72:@6411.4]
  assign _T_10909 = {_T_9864,_T_9863,_T_9862,_T_9861,_T_9860,_T_9859,_T_9858,_T_9857,_T_10901}; // @[Mux.scala 19:72:@6419.4]
  assign _T_10911 = _T_4523 ? _T_10909 : 16'h0; // @[Mux.scala 19:72:@6420.4]
  assign _T_10918 = {_T_9927,_T_9926,_T_9925,_T_9924,_T_9923,_T_9938,_T_9937,_T_9936}; // @[Mux.scala 19:72:@6427.4]
  assign _T_10926 = {_T_9935,_T_9934,_T_9933,_T_9932,_T_9931,_T_9930,_T_9929,_T_9928,_T_10918}; // @[Mux.scala 19:72:@6435.4]
  assign _T_10928 = _T_4524 ? _T_10926 : 16'h0; // @[Mux.scala 19:72:@6436.4]
  assign _T_10935 = {_T_9998,_T_9997,_T_9996,_T_9995,_T_10010,_T_10009,_T_10008,_T_10007}; // @[Mux.scala 19:72:@6443.4]
  assign _T_10943 = {_T_10006,_T_10005,_T_10004,_T_10003,_T_10002,_T_10001,_T_10000,_T_9999,_T_10935}; // @[Mux.scala 19:72:@6451.4]
  assign _T_10945 = _T_4525 ? _T_10943 : 16'h0; // @[Mux.scala 19:72:@6452.4]
  assign _T_10952 = {_T_10069,_T_10068,_T_10067,_T_10082,_T_10081,_T_10080,_T_10079,_T_10078}; // @[Mux.scala 19:72:@6459.4]
  assign _T_10960 = {_T_10077,_T_10076,_T_10075,_T_10074,_T_10073,_T_10072,_T_10071,_T_10070,_T_10952}; // @[Mux.scala 19:72:@6467.4]
  assign _T_10962 = _T_4526 ? _T_10960 : 16'h0; // @[Mux.scala 19:72:@6468.4]
  assign _T_10969 = {_T_10140,_T_10139,_T_10154,_T_10153,_T_10152,_T_10151,_T_10150,_T_10149}; // @[Mux.scala 19:72:@6475.4]
  assign _T_10977 = {_T_10148,_T_10147,_T_10146,_T_10145,_T_10144,_T_10143,_T_10142,_T_10141,_T_10969}; // @[Mux.scala 19:72:@6483.4]
  assign _T_10979 = _T_4527 ? _T_10977 : 16'h0; // @[Mux.scala 19:72:@6484.4]
  assign _T_10986 = {_T_10211,_T_10226,_T_10225,_T_10224,_T_10223,_T_10222,_T_10221,_T_10220}; // @[Mux.scala 19:72:@6491.4]
  assign _T_10994 = {_T_10219,_T_10218,_T_10217,_T_10216,_T_10215,_T_10214,_T_10213,_T_10212,_T_10986}; // @[Mux.scala 19:72:@6499.4]
  assign _T_10996 = _T_4528 ? _T_10994 : 16'h0; // @[Mux.scala 19:72:@6500.4]
  assign _T_11003 = {_T_10298,_T_10297,_T_10296,_T_10295,_T_10294,_T_10293,_T_10292,_T_10291}; // @[Mux.scala 19:72:@6507.4]
  assign _T_11011 = {_T_10290,_T_10289,_T_10288,_T_10287,_T_10286,_T_10285,_T_10284,_T_10283,_T_11003}; // @[Mux.scala 19:72:@6515.4]
  assign _T_11013 = _T_4529 ? _T_11011 : 16'h0; // @[Mux.scala 19:72:@6516.4]
  assign _T_11020 = {_T_10369,_T_10368,_T_10367,_T_10366,_T_10365,_T_10364,_T_10363,_T_10362}; // @[Mux.scala 19:72:@6523.4]
  assign _T_11028 = {_T_10361,_T_10360,_T_10359,_T_10358,_T_10357,_T_10356,_T_10355,_T_10370,_T_11020}; // @[Mux.scala 19:72:@6531.4]
  assign _T_11030 = _T_4530 ? _T_11028 : 16'h0; // @[Mux.scala 19:72:@6532.4]
  assign _T_11037 = {_T_10440,_T_10439,_T_10438,_T_10437,_T_10436,_T_10435,_T_10434,_T_10433}; // @[Mux.scala 19:72:@6539.4]
  assign _T_11045 = {_T_10432,_T_10431,_T_10430,_T_10429,_T_10428,_T_10427,_T_10442,_T_10441,_T_11037}; // @[Mux.scala 19:72:@6547.4]
  assign _T_11047 = _T_4531 ? _T_11045 : 16'h0; // @[Mux.scala 19:72:@6548.4]
  assign _T_11054 = {_T_10511,_T_10510,_T_10509,_T_10508,_T_10507,_T_10506,_T_10505,_T_10504}; // @[Mux.scala 19:72:@6555.4]
  assign _T_11062 = {_T_10503,_T_10502,_T_10501,_T_10500,_T_10499,_T_10514,_T_10513,_T_10512,_T_11054}; // @[Mux.scala 19:72:@6563.4]
  assign _T_11064 = _T_4532 ? _T_11062 : 16'h0; // @[Mux.scala 19:72:@6564.4]
  assign _T_11071 = {_T_10582,_T_10581,_T_10580,_T_10579,_T_10578,_T_10577,_T_10576,_T_10575}; // @[Mux.scala 19:72:@6571.4]
  assign _T_11079 = {_T_10574,_T_10573,_T_10572,_T_10571,_T_10586,_T_10585,_T_10584,_T_10583,_T_11071}; // @[Mux.scala 19:72:@6579.4]
  assign _T_11081 = _T_4533 ? _T_11079 : 16'h0; // @[Mux.scala 19:72:@6580.4]
  assign _T_11088 = {_T_10653,_T_10652,_T_10651,_T_10650,_T_10649,_T_10648,_T_10647,_T_10646}; // @[Mux.scala 19:72:@6587.4]
  assign _T_11096 = {_T_10645,_T_10644,_T_10643,_T_10658,_T_10657,_T_10656,_T_10655,_T_10654,_T_11088}; // @[Mux.scala 19:72:@6595.4]
  assign _T_11098 = _T_4534 ? _T_11096 : 16'h0; // @[Mux.scala 19:72:@6596.4]
  assign _T_11105 = {_T_10724,_T_10723,_T_10722,_T_10721,_T_10720,_T_10719,_T_10718,_T_10717}; // @[Mux.scala 19:72:@6603.4]
  assign _T_11113 = {_T_10716,_T_10715,_T_10730,_T_10729,_T_10728,_T_10727,_T_10726,_T_10725,_T_11105}; // @[Mux.scala 19:72:@6611.4]
  assign _T_11115 = _T_4535 ? _T_11113 : 16'h0; // @[Mux.scala 19:72:@6612.4]
  assign _T_11122 = {_T_10795,_T_10794,_T_10793,_T_10792,_T_10791,_T_10790,_T_10789,_T_10788}; // @[Mux.scala 19:72:@6619.4]
  assign _T_11130 = {_T_10787,_T_10802,_T_10801,_T_10800,_T_10799,_T_10798,_T_10797,_T_10796,_T_11122}; // @[Mux.scala 19:72:@6627.4]
  assign _T_11132 = _T_4536 ? _T_11130 : 16'h0; // @[Mux.scala 19:72:@6628.4]
  assign _T_11133 = _T_10877 | _T_10894; // @[Mux.scala 19:72:@6629.4]
  assign _T_11134 = _T_11133 | _T_10911; // @[Mux.scala 19:72:@6630.4]
  assign _T_11135 = _T_11134 | _T_10928; // @[Mux.scala 19:72:@6631.4]
  assign _T_11136 = _T_11135 | _T_10945; // @[Mux.scala 19:72:@6632.4]
  assign _T_11137 = _T_11136 | _T_10962; // @[Mux.scala 19:72:@6633.4]
  assign _T_11138 = _T_11137 | _T_10979; // @[Mux.scala 19:72:@6634.4]
  assign _T_11139 = _T_11138 | _T_10996; // @[Mux.scala 19:72:@6635.4]
  assign _T_11140 = _T_11139 | _T_11013; // @[Mux.scala 19:72:@6636.4]
  assign _T_11141 = _T_11140 | _T_11030; // @[Mux.scala 19:72:@6637.4]
  assign _T_11142 = _T_11141 | _T_11047; // @[Mux.scala 19:72:@6638.4]
  assign _T_11143 = _T_11142 | _T_11064; // @[Mux.scala 19:72:@6639.4]
  assign _T_11144 = _T_11143 | _T_11081; // @[Mux.scala 19:72:@6640.4]
  assign _T_11145 = _T_11144 | _T_11098; // @[Mux.scala 19:72:@6641.4]
  assign _T_11146 = _T_11145 | _T_11115; // @[Mux.scala 19:72:@6642.4]
  assign _T_11147 = _T_11146 | _T_11132; // @[Mux.scala 19:72:@6643.4]
  assign inputDataPriorityPorts_1_0 = _T_11147[0]; // @[Mux.scala 19:72:@6647.4]
  assign inputDataPriorityPorts_1_1 = _T_11147[1]; // @[Mux.scala 19:72:@6649.4]
  assign inputDataPriorityPorts_1_2 = _T_11147[2]; // @[Mux.scala 19:72:@6651.4]
  assign inputDataPriorityPorts_1_3 = _T_11147[3]; // @[Mux.scala 19:72:@6653.4]
  assign inputDataPriorityPorts_1_4 = _T_11147[4]; // @[Mux.scala 19:72:@6655.4]
  assign inputDataPriorityPorts_1_5 = _T_11147[5]; // @[Mux.scala 19:72:@6657.4]
  assign inputDataPriorityPorts_1_6 = _T_11147[6]; // @[Mux.scala 19:72:@6659.4]
  assign inputDataPriorityPorts_1_7 = _T_11147[7]; // @[Mux.scala 19:72:@6661.4]
  assign inputDataPriorityPorts_1_8 = _T_11147[8]; // @[Mux.scala 19:72:@6663.4]
  assign inputDataPriorityPorts_1_9 = _T_11147[9]; // @[Mux.scala 19:72:@6665.4]
  assign inputDataPriorityPorts_1_10 = _T_11147[10]; // @[Mux.scala 19:72:@6667.4]
  assign inputDataPriorityPorts_1_11 = _T_11147[11]; // @[Mux.scala 19:72:@6669.4]
  assign inputDataPriorityPorts_1_12 = _T_11147[12]; // @[Mux.scala 19:72:@6671.4]
  assign inputDataPriorityPorts_1_13 = _T_11147[13]; // @[Mux.scala 19:72:@6673.4]
  assign inputDataPriorityPorts_1_14 = _T_11147[14]; // @[Mux.scala 19:72:@6675.4]
  assign inputDataPriorityPorts_1_15 = _T_11147[15]; // @[Mux.scala 19:72:@6677.4]
  assign _T_11293 = inputAddrPriorityPorts_0_0 & _T_4378; // @[StoreQueue.scala 209:52:@6701.6]
  assign _T_11294 = _T_11293 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6702.6]
  assign _T_11297 = inputAddrPriorityPorts_1_0 & _T_4378; // @[StoreQueue.scala 209:52:@6704.6]
  assign _T_11298 = _T_11297 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6705.6]
  assign _T_11309 = _T_11294 | _T_11298; // @[StoreQueue.scala 210:30:@6710.6]
  assign _T_11310 = {_T_11298,_T_11294}; // @[OneHot.scala 18:45:@6712.8]
  assign _T_11311 = _T_11310[1]; // @[CircuitMath.scala 30:8:@6713.8]
  assign _GEN_993 = _T_11311 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6714.8]
  assign _GEN_994 = _T_11309 ? _GEN_993 : addrQ_0; // @[StoreQueue.scala 210:40:@6711.6]
  assign _GEN_995 = _T_11309 ? 1'h1 : addrKnown_0; // @[StoreQueue.scala 210:40:@6711.6]
  assign _T_11316 = inputDataPriorityPorts_0_0 & _T_4448; // @[StoreQueue.scala 215:52:@6718.6]
  assign _T_11317 = _T_11316 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6719.6]
  assign _T_11320 = inputDataPriorityPorts_1_0 & _T_4448; // @[StoreQueue.scala 215:52:@6721.6]
  assign _T_11321 = _T_11320 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6722.6]
  assign _T_11332 = _T_11317 | _T_11321; // @[StoreQueue.scala 216:30:@6727.6]
  assign _T_11333 = {_T_11321,_T_11317}; // @[OneHot.scala 18:45:@6729.8]
  assign _T_11334 = _T_11333[1]; // @[CircuitMath.scala 30:8:@6730.8]
  assign _GEN_997 = _T_11334 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6731.8]
  assign _GEN_998 = _T_11332 ? _GEN_997 : dataQ_0; // @[StoreQueue.scala 216:40:@6728.6]
  assign _GEN_999 = _T_11332 ? 1'h1 : dataKnown_0; // @[StoreQueue.scala 216:40:@6728.6]
  assign _GEN_1000 = initBits_0 ? 1'h0 : _GEN_995; // @[StoreQueue.scala 204:35:@6695.4]
  assign _GEN_1001 = initBits_0 ? 1'h0 : _GEN_999; // @[StoreQueue.scala 204:35:@6695.4]
  assign _GEN_1002 = initBits_0 ? addrQ_0 : _GEN_994; // @[StoreQueue.scala 204:35:@6695.4]
  assign _GEN_1003 = initBits_0 ? dataQ_0 : _GEN_998; // @[StoreQueue.scala 204:35:@6695.4]
  assign _T_11341 = inputAddrPriorityPorts_0_1 & _T_4381; // @[StoreQueue.scala 209:52:@6741.6]
  assign _T_11342 = _T_11341 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6742.6]
  assign _T_11345 = inputAddrPriorityPorts_1_1 & _T_4381; // @[StoreQueue.scala 209:52:@6744.6]
  assign _T_11346 = _T_11345 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6745.6]
  assign _T_11357 = _T_11342 | _T_11346; // @[StoreQueue.scala 210:30:@6750.6]
  assign _T_11358 = {_T_11346,_T_11342}; // @[OneHot.scala 18:45:@6752.8]
  assign _T_11359 = _T_11358[1]; // @[CircuitMath.scala 30:8:@6753.8]
  assign _GEN_1005 = _T_11359 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6754.8]
  assign _GEN_1006 = _T_11357 ? _GEN_1005 : addrQ_1; // @[StoreQueue.scala 210:40:@6751.6]
  assign _GEN_1007 = _T_11357 ? 1'h1 : addrKnown_1; // @[StoreQueue.scala 210:40:@6751.6]
  assign _T_11364 = inputDataPriorityPorts_0_1 & _T_4451; // @[StoreQueue.scala 215:52:@6758.6]
  assign _T_11365 = _T_11364 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6759.6]
  assign _T_11368 = inputDataPriorityPorts_1_1 & _T_4451; // @[StoreQueue.scala 215:52:@6761.6]
  assign _T_11369 = _T_11368 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6762.6]
  assign _T_11380 = _T_11365 | _T_11369; // @[StoreQueue.scala 216:30:@6767.6]
  assign _T_11381 = {_T_11369,_T_11365}; // @[OneHot.scala 18:45:@6769.8]
  assign _T_11382 = _T_11381[1]; // @[CircuitMath.scala 30:8:@6770.8]
  assign _GEN_1009 = _T_11382 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6771.8]
  assign _GEN_1010 = _T_11380 ? _GEN_1009 : dataQ_1; // @[StoreQueue.scala 216:40:@6768.6]
  assign _GEN_1011 = _T_11380 ? 1'h1 : dataKnown_1; // @[StoreQueue.scala 216:40:@6768.6]
  assign _GEN_1012 = initBits_1 ? 1'h0 : _GEN_1007; // @[StoreQueue.scala 204:35:@6735.4]
  assign _GEN_1013 = initBits_1 ? 1'h0 : _GEN_1011; // @[StoreQueue.scala 204:35:@6735.4]
  assign _GEN_1014 = initBits_1 ? addrQ_1 : _GEN_1006; // @[StoreQueue.scala 204:35:@6735.4]
  assign _GEN_1015 = initBits_1 ? dataQ_1 : _GEN_1010; // @[StoreQueue.scala 204:35:@6735.4]
  assign _T_11389 = inputAddrPriorityPorts_0_2 & _T_4384; // @[StoreQueue.scala 209:52:@6781.6]
  assign _T_11390 = _T_11389 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6782.6]
  assign _T_11393 = inputAddrPriorityPorts_1_2 & _T_4384; // @[StoreQueue.scala 209:52:@6784.6]
  assign _T_11394 = _T_11393 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6785.6]
  assign _T_11405 = _T_11390 | _T_11394; // @[StoreQueue.scala 210:30:@6790.6]
  assign _T_11406 = {_T_11394,_T_11390}; // @[OneHot.scala 18:45:@6792.8]
  assign _T_11407 = _T_11406[1]; // @[CircuitMath.scala 30:8:@6793.8]
  assign _GEN_1017 = _T_11407 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6794.8]
  assign _GEN_1018 = _T_11405 ? _GEN_1017 : addrQ_2; // @[StoreQueue.scala 210:40:@6791.6]
  assign _GEN_1019 = _T_11405 ? 1'h1 : addrKnown_2; // @[StoreQueue.scala 210:40:@6791.6]
  assign _T_11412 = inputDataPriorityPorts_0_2 & _T_4454; // @[StoreQueue.scala 215:52:@6798.6]
  assign _T_11413 = _T_11412 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6799.6]
  assign _T_11416 = inputDataPriorityPorts_1_2 & _T_4454; // @[StoreQueue.scala 215:52:@6801.6]
  assign _T_11417 = _T_11416 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6802.6]
  assign _T_11428 = _T_11413 | _T_11417; // @[StoreQueue.scala 216:30:@6807.6]
  assign _T_11429 = {_T_11417,_T_11413}; // @[OneHot.scala 18:45:@6809.8]
  assign _T_11430 = _T_11429[1]; // @[CircuitMath.scala 30:8:@6810.8]
  assign _GEN_1021 = _T_11430 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6811.8]
  assign _GEN_1022 = _T_11428 ? _GEN_1021 : dataQ_2; // @[StoreQueue.scala 216:40:@6808.6]
  assign _GEN_1023 = _T_11428 ? 1'h1 : dataKnown_2; // @[StoreQueue.scala 216:40:@6808.6]
  assign _GEN_1024 = initBits_2 ? 1'h0 : _GEN_1019; // @[StoreQueue.scala 204:35:@6775.4]
  assign _GEN_1025 = initBits_2 ? 1'h0 : _GEN_1023; // @[StoreQueue.scala 204:35:@6775.4]
  assign _GEN_1026 = initBits_2 ? addrQ_2 : _GEN_1018; // @[StoreQueue.scala 204:35:@6775.4]
  assign _GEN_1027 = initBits_2 ? dataQ_2 : _GEN_1022; // @[StoreQueue.scala 204:35:@6775.4]
  assign _T_11437 = inputAddrPriorityPorts_0_3 & _T_4387; // @[StoreQueue.scala 209:52:@6821.6]
  assign _T_11438 = _T_11437 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6822.6]
  assign _T_11441 = inputAddrPriorityPorts_1_3 & _T_4387; // @[StoreQueue.scala 209:52:@6824.6]
  assign _T_11442 = _T_11441 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6825.6]
  assign _T_11453 = _T_11438 | _T_11442; // @[StoreQueue.scala 210:30:@6830.6]
  assign _T_11454 = {_T_11442,_T_11438}; // @[OneHot.scala 18:45:@6832.8]
  assign _T_11455 = _T_11454[1]; // @[CircuitMath.scala 30:8:@6833.8]
  assign _GEN_1029 = _T_11455 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6834.8]
  assign _GEN_1030 = _T_11453 ? _GEN_1029 : addrQ_3; // @[StoreQueue.scala 210:40:@6831.6]
  assign _GEN_1031 = _T_11453 ? 1'h1 : addrKnown_3; // @[StoreQueue.scala 210:40:@6831.6]
  assign _T_11460 = inputDataPriorityPorts_0_3 & _T_4457; // @[StoreQueue.scala 215:52:@6838.6]
  assign _T_11461 = _T_11460 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6839.6]
  assign _T_11464 = inputDataPriorityPorts_1_3 & _T_4457; // @[StoreQueue.scala 215:52:@6841.6]
  assign _T_11465 = _T_11464 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6842.6]
  assign _T_11476 = _T_11461 | _T_11465; // @[StoreQueue.scala 216:30:@6847.6]
  assign _T_11477 = {_T_11465,_T_11461}; // @[OneHot.scala 18:45:@6849.8]
  assign _T_11478 = _T_11477[1]; // @[CircuitMath.scala 30:8:@6850.8]
  assign _GEN_1033 = _T_11478 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6851.8]
  assign _GEN_1034 = _T_11476 ? _GEN_1033 : dataQ_3; // @[StoreQueue.scala 216:40:@6848.6]
  assign _GEN_1035 = _T_11476 ? 1'h1 : dataKnown_3; // @[StoreQueue.scala 216:40:@6848.6]
  assign _GEN_1036 = initBits_3 ? 1'h0 : _GEN_1031; // @[StoreQueue.scala 204:35:@6815.4]
  assign _GEN_1037 = initBits_3 ? 1'h0 : _GEN_1035; // @[StoreQueue.scala 204:35:@6815.4]
  assign _GEN_1038 = initBits_3 ? addrQ_3 : _GEN_1030; // @[StoreQueue.scala 204:35:@6815.4]
  assign _GEN_1039 = initBits_3 ? dataQ_3 : _GEN_1034; // @[StoreQueue.scala 204:35:@6815.4]
  assign _T_11485 = inputAddrPriorityPorts_0_4 & _T_4390; // @[StoreQueue.scala 209:52:@6861.6]
  assign _T_11486 = _T_11485 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6862.6]
  assign _T_11489 = inputAddrPriorityPorts_1_4 & _T_4390; // @[StoreQueue.scala 209:52:@6864.6]
  assign _T_11490 = _T_11489 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6865.6]
  assign _T_11501 = _T_11486 | _T_11490; // @[StoreQueue.scala 210:30:@6870.6]
  assign _T_11502 = {_T_11490,_T_11486}; // @[OneHot.scala 18:45:@6872.8]
  assign _T_11503 = _T_11502[1]; // @[CircuitMath.scala 30:8:@6873.8]
  assign _GEN_1041 = _T_11503 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6874.8]
  assign _GEN_1042 = _T_11501 ? _GEN_1041 : addrQ_4; // @[StoreQueue.scala 210:40:@6871.6]
  assign _GEN_1043 = _T_11501 ? 1'h1 : addrKnown_4; // @[StoreQueue.scala 210:40:@6871.6]
  assign _T_11508 = inputDataPriorityPorts_0_4 & _T_4460; // @[StoreQueue.scala 215:52:@6878.6]
  assign _T_11509 = _T_11508 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6879.6]
  assign _T_11512 = inputDataPriorityPorts_1_4 & _T_4460; // @[StoreQueue.scala 215:52:@6881.6]
  assign _T_11513 = _T_11512 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6882.6]
  assign _T_11524 = _T_11509 | _T_11513; // @[StoreQueue.scala 216:30:@6887.6]
  assign _T_11525 = {_T_11513,_T_11509}; // @[OneHot.scala 18:45:@6889.8]
  assign _T_11526 = _T_11525[1]; // @[CircuitMath.scala 30:8:@6890.8]
  assign _GEN_1045 = _T_11526 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6891.8]
  assign _GEN_1046 = _T_11524 ? _GEN_1045 : dataQ_4; // @[StoreQueue.scala 216:40:@6888.6]
  assign _GEN_1047 = _T_11524 ? 1'h1 : dataKnown_4; // @[StoreQueue.scala 216:40:@6888.6]
  assign _GEN_1048 = initBits_4 ? 1'h0 : _GEN_1043; // @[StoreQueue.scala 204:35:@6855.4]
  assign _GEN_1049 = initBits_4 ? 1'h0 : _GEN_1047; // @[StoreQueue.scala 204:35:@6855.4]
  assign _GEN_1050 = initBits_4 ? addrQ_4 : _GEN_1042; // @[StoreQueue.scala 204:35:@6855.4]
  assign _GEN_1051 = initBits_4 ? dataQ_4 : _GEN_1046; // @[StoreQueue.scala 204:35:@6855.4]
  assign _T_11533 = inputAddrPriorityPorts_0_5 & _T_4393; // @[StoreQueue.scala 209:52:@6901.6]
  assign _T_11534 = _T_11533 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6902.6]
  assign _T_11537 = inputAddrPriorityPorts_1_5 & _T_4393; // @[StoreQueue.scala 209:52:@6904.6]
  assign _T_11538 = _T_11537 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6905.6]
  assign _T_11549 = _T_11534 | _T_11538; // @[StoreQueue.scala 210:30:@6910.6]
  assign _T_11550 = {_T_11538,_T_11534}; // @[OneHot.scala 18:45:@6912.8]
  assign _T_11551 = _T_11550[1]; // @[CircuitMath.scala 30:8:@6913.8]
  assign _GEN_1053 = _T_11551 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6914.8]
  assign _GEN_1054 = _T_11549 ? _GEN_1053 : addrQ_5; // @[StoreQueue.scala 210:40:@6911.6]
  assign _GEN_1055 = _T_11549 ? 1'h1 : addrKnown_5; // @[StoreQueue.scala 210:40:@6911.6]
  assign _T_11556 = inputDataPriorityPorts_0_5 & _T_4463; // @[StoreQueue.scala 215:52:@6918.6]
  assign _T_11557 = _T_11556 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6919.6]
  assign _T_11560 = inputDataPriorityPorts_1_5 & _T_4463; // @[StoreQueue.scala 215:52:@6921.6]
  assign _T_11561 = _T_11560 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6922.6]
  assign _T_11572 = _T_11557 | _T_11561; // @[StoreQueue.scala 216:30:@6927.6]
  assign _T_11573 = {_T_11561,_T_11557}; // @[OneHot.scala 18:45:@6929.8]
  assign _T_11574 = _T_11573[1]; // @[CircuitMath.scala 30:8:@6930.8]
  assign _GEN_1057 = _T_11574 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6931.8]
  assign _GEN_1058 = _T_11572 ? _GEN_1057 : dataQ_5; // @[StoreQueue.scala 216:40:@6928.6]
  assign _GEN_1059 = _T_11572 ? 1'h1 : dataKnown_5; // @[StoreQueue.scala 216:40:@6928.6]
  assign _GEN_1060 = initBits_5 ? 1'h0 : _GEN_1055; // @[StoreQueue.scala 204:35:@6895.4]
  assign _GEN_1061 = initBits_5 ? 1'h0 : _GEN_1059; // @[StoreQueue.scala 204:35:@6895.4]
  assign _GEN_1062 = initBits_5 ? addrQ_5 : _GEN_1054; // @[StoreQueue.scala 204:35:@6895.4]
  assign _GEN_1063 = initBits_5 ? dataQ_5 : _GEN_1058; // @[StoreQueue.scala 204:35:@6895.4]
  assign _T_11581 = inputAddrPriorityPorts_0_6 & _T_4396; // @[StoreQueue.scala 209:52:@6941.6]
  assign _T_11582 = _T_11581 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6942.6]
  assign _T_11585 = inputAddrPriorityPorts_1_6 & _T_4396; // @[StoreQueue.scala 209:52:@6944.6]
  assign _T_11586 = _T_11585 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6945.6]
  assign _T_11597 = _T_11582 | _T_11586; // @[StoreQueue.scala 210:30:@6950.6]
  assign _T_11598 = {_T_11586,_T_11582}; // @[OneHot.scala 18:45:@6952.8]
  assign _T_11599 = _T_11598[1]; // @[CircuitMath.scala 30:8:@6953.8]
  assign _GEN_1065 = _T_11599 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6954.8]
  assign _GEN_1066 = _T_11597 ? _GEN_1065 : addrQ_6; // @[StoreQueue.scala 210:40:@6951.6]
  assign _GEN_1067 = _T_11597 ? 1'h1 : addrKnown_6; // @[StoreQueue.scala 210:40:@6951.6]
  assign _T_11604 = inputDataPriorityPorts_0_6 & _T_4466; // @[StoreQueue.scala 215:52:@6958.6]
  assign _T_11605 = _T_11604 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6959.6]
  assign _T_11608 = inputDataPriorityPorts_1_6 & _T_4466; // @[StoreQueue.scala 215:52:@6961.6]
  assign _T_11609 = _T_11608 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@6962.6]
  assign _T_11620 = _T_11605 | _T_11609; // @[StoreQueue.scala 216:30:@6967.6]
  assign _T_11621 = {_T_11609,_T_11605}; // @[OneHot.scala 18:45:@6969.8]
  assign _T_11622 = _T_11621[1]; // @[CircuitMath.scala 30:8:@6970.8]
  assign _GEN_1069 = _T_11622 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@6971.8]
  assign _GEN_1070 = _T_11620 ? _GEN_1069 : dataQ_6; // @[StoreQueue.scala 216:40:@6968.6]
  assign _GEN_1071 = _T_11620 ? 1'h1 : dataKnown_6; // @[StoreQueue.scala 216:40:@6968.6]
  assign _GEN_1072 = initBits_6 ? 1'h0 : _GEN_1067; // @[StoreQueue.scala 204:35:@6935.4]
  assign _GEN_1073 = initBits_6 ? 1'h0 : _GEN_1071; // @[StoreQueue.scala 204:35:@6935.4]
  assign _GEN_1074 = initBits_6 ? addrQ_6 : _GEN_1066; // @[StoreQueue.scala 204:35:@6935.4]
  assign _GEN_1075 = initBits_6 ? dataQ_6 : _GEN_1070; // @[StoreQueue.scala 204:35:@6935.4]
  assign _T_11629 = inputAddrPriorityPorts_0_7 & _T_4399; // @[StoreQueue.scala 209:52:@6981.6]
  assign _T_11630 = _T_11629 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@6982.6]
  assign _T_11633 = inputAddrPriorityPorts_1_7 & _T_4399; // @[StoreQueue.scala 209:52:@6984.6]
  assign _T_11634 = _T_11633 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@6985.6]
  assign _T_11645 = _T_11630 | _T_11634; // @[StoreQueue.scala 210:30:@6990.6]
  assign _T_11646 = {_T_11634,_T_11630}; // @[OneHot.scala 18:45:@6992.8]
  assign _T_11647 = _T_11646[1]; // @[CircuitMath.scala 30:8:@6993.8]
  assign _GEN_1077 = _T_11647 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@6994.8]
  assign _GEN_1078 = _T_11645 ? _GEN_1077 : addrQ_7; // @[StoreQueue.scala 210:40:@6991.6]
  assign _GEN_1079 = _T_11645 ? 1'h1 : addrKnown_7; // @[StoreQueue.scala 210:40:@6991.6]
  assign _T_11652 = inputDataPriorityPorts_0_7 & _T_4469; // @[StoreQueue.scala 215:52:@6998.6]
  assign _T_11653 = _T_11652 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@6999.6]
  assign _T_11656 = inputDataPriorityPorts_1_7 & _T_4469; // @[StoreQueue.scala 215:52:@7001.6]
  assign _T_11657 = _T_11656 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7002.6]
  assign _T_11668 = _T_11653 | _T_11657; // @[StoreQueue.scala 216:30:@7007.6]
  assign _T_11669 = {_T_11657,_T_11653}; // @[OneHot.scala 18:45:@7009.8]
  assign _T_11670 = _T_11669[1]; // @[CircuitMath.scala 30:8:@7010.8]
  assign _GEN_1081 = _T_11670 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7011.8]
  assign _GEN_1082 = _T_11668 ? _GEN_1081 : dataQ_7; // @[StoreQueue.scala 216:40:@7008.6]
  assign _GEN_1083 = _T_11668 ? 1'h1 : dataKnown_7; // @[StoreQueue.scala 216:40:@7008.6]
  assign _GEN_1084 = initBits_7 ? 1'h0 : _GEN_1079; // @[StoreQueue.scala 204:35:@6975.4]
  assign _GEN_1085 = initBits_7 ? 1'h0 : _GEN_1083; // @[StoreQueue.scala 204:35:@6975.4]
  assign _GEN_1086 = initBits_7 ? addrQ_7 : _GEN_1078; // @[StoreQueue.scala 204:35:@6975.4]
  assign _GEN_1087 = initBits_7 ? dataQ_7 : _GEN_1082; // @[StoreQueue.scala 204:35:@6975.4]
  assign _T_11677 = inputAddrPriorityPorts_0_8 & _T_4402; // @[StoreQueue.scala 209:52:@7021.6]
  assign _T_11678 = _T_11677 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7022.6]
  assign _T_11681 = inputAddrPriorityPorts_1_8 & _T_4402; // @[StoreQueue.scala 209:52:@7024.6]
  assign _T_11682 = _T_11681 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7025.6]
  assign _T_11693 = _T_11678 | _T_11682; // @[StoreQueue.scala 210:30:@7030.6]
  assign _T_11694 = {_T_11682,_T_11678}; // @[OneHot.scala 18:45:@7032.8]
  assign _T_11695 = _T_11694[1]; // @[CircuitMath.scala 30:8:@7033.8]
  assign _GEN_1089 = _T_11695 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7034.8]
  assign _GEN_1090 = _T_11693 ? _GEN_1089 : addrQ_8; // @[StoreQueue.scala 210:40:@7031.6]
  assign _GEN_1091 = _T_11693 ? 1'h1 : addrKnown_8; // @[StoreQueue.scala 210:40:@7031.6]
  assign _T_11700 = inputDataPriorityPorts_0_8 & _T_4472; // @[StoreQueue.scala 215:52:@7038.6]
  assign _T_11701 = _T_11700 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7039.6]
  assign _T_11704 = inputDataPriorityPorts_1_8 & _T_4472; // @[StoreQueue.scala 215:52:@7041.6]
  assign _T_11705 = _T_11704 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7042.6]
  assign _T_11716 = _T_11701 | _T_11705; // @[StoreQueue.scala 216:30:@7047.6]
  assign _T_11717 = {_T_11705,_T_11701}; // @[OneHot.scala 18:45:@7049.8]
  assign _T_11718 = _T_11717[1]; // @[CircuitMath.scala 30:8:@7050.8]
  assign _GEN_1093 = _T_11718 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7051.8]
  assign _GEN_1094 = _T_11716 ? _GEN_1093 : dataQ_8; // @[StoreQueue.scala 216:40:@7048.6]
  assign _GEN_1095 = _T_11716 ? 1'h1 : dataKnown_8; // @[StoreQueue.scala 216:40:@7048.6]
  assign _GEN_1096 = initBits_8 ? 1'h0 : _GEN_1091; // @[StoreQueue.scala 204:35:@7015.4]
  assign _GEN_1097 = initBits_8 ? 1'h0 : _GEN_1095; // @[StoreQueue.scala 204:35:@7015.4]
  assign _GEN_1098 = initBits_8 ? addrQ_8 : _GEN_1090; // @[StoreQueue.scala 204:35:@7015.4]
  assign _GEN_1099 = initBits_8 ? dataQ_8 : _GEN_1094; // @[StoreQueue.scala 204:35:@7015.4]
  assign _T_11725 = inputAddrPriorityPorts_0_9 & _T_4405; // @[StoreQueue.scala 209:52:@7061.6]
  assign _T_11726 = _T_11725 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7062.6]
  assign _T_11729 = inputAddrPriorityPorts_1_9 & _T_4405; // @[StoreQueue.scala 209:52:@7064.6]
  assign _T_11730 = _T_11729 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7065.6]
  assign _T_11741 = _T_11726 | _T_11730; // @[StoreQueue.scala 210:30:@7070.6]
  assign _T_11742 = {_T_11730,_T_11726}; // @[OneHot.scala 18:45:@7072.8]
  assign _T_11743 = _T_11742[1]; // @[CircuitMath.scala 30:8:@7073.8]
  assign _GEN_1101 = _T_11743 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7074.8]
  assign _GEN_1102 = _T_11741 ? _GEN_1101 : addrQ_9; // @[StoreQueue.scala 210:40:@7071.6]
  assign _GEN_1103 = _T_11741 ? 1'h1 : addrKnown_9; // @[StoreQueue.scala 210:40:@7071.6]
  assign _T_11748 = inputDataPriorityPorts_0_9 & _T_4475; // @[StoreQueue.scala 215:52:@7078.6]
  assign _T_11749 = _T_11748 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7079.6]
  assign _T_11752 = inputDataPriorityPorts_1_9 & _T_4475; // @[StoreQueue.scala 215:52:@7081.6]
  assign _T_11753 = _T_11752 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7082.6]
  assign _T_11764 = _T_11749 | _T_11753; // @[StoreQueue.scala 216:30:@7087.6]
  assign _T_11765 = {_T_11753,_T_11749}; // @[OneHot.scala 18:45:@7089.8]
  assign _T_11766 = _T_11765[1]; // @[CircuitMath.scala 30:8:@7090.8]
  assign _GEN_1105 = _T_11766 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7091.8]
  assign _GEN_1106 = _T_11764 ? _GEN_1105 : dataQ_9; // @[StoreQueue.scala 216:40:@7088.6]
  assign _GEN_1107 = _T_11764 ? 1'h1 : dataKnown_9; // @[StoreQueue.scala 216:40:@7088.6]
  assign _GEN_1108 = initBits_9 ? 1'h0 : _GEN_1103; // @[StoreQueue.scala 204:35:@7055.4]
  assign _GEN_1109 = initBits_9 ? 1'h0 : _GEN_1107; // @[StoreQueue.scala 204:35:@7055.4]
  assign _GEN_1110 = initBits_9 ? addrQ_9 : _GEN_1102; // @[StoreQueue.scala 204:35:@7055.4]
  assign _GEN_1111 = initBits_9 ? dataQ_9 : _GEN_1106; // @[StoreQueue.scala 204:35:@7055.4]
  assign _T_11773 = inputAddrPriorityPorts_0_10 & _T_4408; // @[StoreQueue.scala 209:52:@7101.6]
  assign _T_11774 = _T_11773 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7102.6]
  assign _T_11777 = inputAddrPriorityPorts_1_10 & _T_4408; // @[StoreQueue.scala 209:52:@7104.6]
  assign _T_11778 = _T_11777 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7105.6]
  assign _T_11789 = _T_11774 | _T_11778; // @[StoreQueue.scala 210:30:@7110.6]
  assign _T_11790 = {_T_11778,_T_11774}; // @[OneHot.scala 18:45:@7112.8]
  assign _T_11791 = _T_11790[1]; // @[CircuitMath.scala 30:8:@7113.8]
  assign _GEN_1113 = _T_11791 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7114.8]
  assign _GEN_1114 = _T_11789 ? _GEN_1113 : addrQ_10; // @[StoreQueue.scala 210:40:@7111.6]
  assign _GEN_1115 = _T_11789 ? 1'h1 : addrKnown_10; // @[StoreQueue.scala 210:40:@7111.6]
  assign _T_11796 = inputDataPriorityPorts_0_10 & _T_4478; // @[StoreQueue.scala 215:52:@7118.6]
  assign _T_11797 = _T_11796 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7119.6]
  assign _T_11800 = inputDataPriorityPorts_1_10 & _T_4478; // @[StoreQueue.scala 215:52:@7121.6]
  assign _T_11801 = _T_11800 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7122.6]
  assign _T_11812 = _T_11797 | _T_11801; // @[StoreQueue.scala 216:30:@7127.6]
  assign _T_11813 = {_T_11801,_T_11797}; // @[OneHot.scala 18:45:@7129.8]
  assign _T_11814 = _T_11813[1]; // @[CircuitMath.scala 30:8:@7130.8]
  assign _GEN_1117 = _T_11814 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7131.8]
  assign _GEN_1118 = _T_11812 ? _GEN_1117 : dataQ_10; // @[StoreQueue.scala 216:40:@7128.6]
  assign _GEN_1119 = _T_11812 ? 1'h1 : dataKnown_10; // @[StoreQueue.scala 216:40:@7128.6]
  assign _GEN_1120 = initBits_10 ? 1'h0 : _GEN_1115; // @[StoreQueue.scala 204:35:@7095.4]
  assign _GEN_1121 = initBits_10 ? 1'h0 : _GEN_1119; // @[StoreQueue.scala 204:35:@7095.4]
  assign _GEN_1122 = initBits_10 ? addrQ_10 : _GEN_1114; // @[StoreQueue.scala 204:35:@7095.4]
  assign _GEN_1123 = initBits_10 ? dataQ_10 : _GEN_1118; // @[StoreQueue.scala 204:35:@7095.4]
  assign _T_11821 = inputAddrPriorityPorts_0_11 & _T_4411; // @[StoreQueue.scala 209:52:@7141.6]
  assign _T_11822 = _T_11821 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7142.6]
  assign _T_11825 = inputAddrPriorityPorts_1_11 & _T_4411; // @[StoreQueue.scala 209:52:@7144.6]
  assign _T_11826 = _T_11825 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7145.6]
  assign _T_11837 = _T_11822 | _T_11826; // @[StoreQueue.scala 210:30:@7150.6]
  assign _T_11838 = {_T_11826,_T_11822}; // @[OneHot.scala 18:45:@7152.8]
  assign _T_11839 = _T_11838[1]; // @[CircuitMath.scala 30:8:@7153.8]
  assign _GEN_1125 = _T_11839 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7154.8]
  assign _GEN_1126 = _T_11837 ? _GEN_1125 : addrQ_11; // @[StoreQueue.scala 210:40:@7151.6]
  assign _GEN_1127 = _T_11837 ? 1'h1 : addrKnown_11; // @[StoreQueue.scala 210:40:@7151.6]
  assign _T_11844 = inputDataPriorityPorts_0_11 & _T_4481; // @[StoreQueue.scala 215:52:@7158.6]
  assign _T_11845 = _T_11844 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7159.6]
  assign _T_11848 = inputDataPriorityPorts_1_11 & _T_4481; // @[StoreQueue.scala 215:52:@7161.6]
  assign _T_11849 = _T_11848 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7162.6]
  assign _T_11860 = _T_11845 | _T_11849; // @[StoreQueue.scala 216:30:@7167.6]
  assign _T_11861 = {_T_11849,_T_11845}; // @[OneHot.scala 18:45:@7169.8]
  assign _T_11862 = _T_11861[1]; // @[CircuitMath.scala 30:8:@7170.8]
  assign _GEN_1129 = _T_11862 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7171.8]
  assign _GEN_1130 = _T_11860 ? _GEN_1129 : dataQ_11; // @[StoreQueue.scala 216:40:@7168.6]
  assign _GEN_1131 = _T_11860 ? 1'h1 : dataKnown_11; // @[StoreQueue.scala 216:40:@7168.6]
  assign _GEN_1132 = initBits_11 ? 1'h0 : _GEN_1127; // @[StoreQueue.scala 204:35:@7135.4]
  assign _GEN_1133 = initBits_11 ? 1'h0 : _GEN_1131; // @[StoreQueue.scala 204:35:@7135.4]
  assign _GEN_1134 = initBits_11 ? addrQ_11 : _GEN_1126; // @[StoreQueue.scala 204:35:@7135.4]
  assign _GEN_1135 = initBits_11 ? dataQ_11 : _GEN_1130; // @[StoreQueue.scala 204:35:@7135.4]
  assign _T_11869 = inputAddrPriorityPorts_0_12 & _T_4414; // @[StoreQueue.scala 209:52:@7181.6]
  assign _T_11870 = _T_11869 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7182.6]
  assign _T_11873 = inputAddrPriorityPorts_1_12 & _T_4414; // @[StoreQueue.scala 209:52:@7184.6]
  assign _T_11874 = _T_11873 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7185.6]
  assign _T_11885 = _T_11870 | _T_11874; // @[StoreQueue.scala 210:30:@7190.6]
  assign _T_11886 = {_T_11874,_T_11870}; // @[OneHot.scala 18:45:@7192.8]
  assign _T_11887 = _T_11886[1]; // @[CircuitMath.scala 30:8:@7193.8]
  assign _GEN_1137 = _T_11887 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7194.8]
  assign _GEN_1138 = _T_11885 ? _GEN_1137 : addrQ_12; // @[StoreQueue.scala 210:40:@7191.6]
  assign _GEN_1139 = _T_11885 ? 1'h1 : addrKnown_12; // @[StoreQueue.scala 210:40:@7191.6]
  assign _T_11892 = inputDataPriorityPorts_0_12 & _T_4484; // @[StoreQueue.scala 215:52:@7198.6]
  assign _T_11893 = _T_11892 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7199.6]
  assign _T_11896 = inputDataPriorityPorts_1_12 & _T_4484; // @[StoreQueue.scala 215:52:@7201.6]
  assign _T_11897 = _T_11896 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7202.6]
  assign _T_11908 = _T_11893 | _T_11897; // @[StoreQueue.scala 216:30:@7207.6]
  assign _T_11909 = {_T_11897,_T_11893}; // @[OneHot.scala 18:45:@7209.8]
  assign _T_11910 = _T_11909[1]; // @[CircuitMath.scala 30:8:@7210.8]
  assign _GEN_1141 = _T_11910 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7211.8]
  assign _GEN_1142 = _T_11908 ? _GEN_1141 : dataQ_12; // @[StoreQueue.scala 216:40:@7208.6]
  assign _GEN_1143 = _T_11908 ? 1'h1 : dataKnown_12; // @[StoreQueue.scala 216:40:@7208.6]
  assign _GEN_1144 = initBits_12 ? 1'h0 : _GEN_1139; // @[StoreQueue.scala 204:35:@7175.4]
  assign _GEN_1145 = initBits_12 ? 1'h0 : _GEN_1143; // @[StoreQueue.scala 204:35:@7175.4]
  assign _GEN_1146 = initBits_12 ? addrQ_12 : _GEN_1138; // @[StoreQueue.scala 204:35:@7175.4]
  assign _GEN_1147 = initBits_12 ? dataQ_12 : _GEN_1142; // @[StoreQueue.scala 204:35:@7175.4]
  assign _T_11917 = inputAddrPriorityPorts_0_13 & _T_4417; // @[StoreQueue.scala 209:52:@7221.6]
  assign _T_11918 = _T_11917 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7222.6]
  assign _T_11921 = inputAddrPriorityPorts_1_13 & _T_4417; // @[StoreQueue.scala 209:52:@7224.6]
  assign _T_11922 = _T_11921 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7225.6]
  assign _T_11933 = _T_11918 | _T_11922; // @[StoreQueue.scala 210:30:@7230.6]
  assign _T_11934 = {_T_11922,_T_11918}; // @[OneHot.scala 18:45:@7232.8]
  assign _T_11935 = _T_11934[1]; // @[CircuitMath.scala 30:8:@7233.8]
  assign _GEN_1149 = _T_11935 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7234.8]
  assign _GEN_1150 = _T_11933 ? _GEN_1149 : addrQ_13; // @[StoreQueue.scala 210:40:@7231.6]
  assign _GEN_1151 = _T_11933 ? 1'h1 : addrKnown_13; // @[StoreQueue.scala 210:40:@7231.6]
  assign _T_11940 = inputDataPriorityPorts_0_13 & _T_4487; // @[StoreQueue.scala 215:52:@7238.6]
  assign _T_11941 = _T_11940 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7239.6]
  assign _T_11944 = inputDataPriorityPorts_1_13 & _T_4487; // @[StoreQueue.scala 215:52:@7241.6]
  assign _T_11945 = _T_11944 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7242.6]
  assign _T_11956 = _T_11941 | _T_11945; // @[StoreQueue.scala 216:30:@7247.6]
  assign _T_11957 = {_T_11945,_T_11941}; // @[OneHot.scala 18:45:@7249.8]
  assign _T_11958 = _T_11957[1]; // @[CircuitMath.scala 30:8:@7250.8]
  assign _GEN_1153 = _T_11958 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7251.8]
  assign _GEN_1154 = _T_11956 ? _GEN_1153 : dataQ_13; // @[StoreQueue.scala 216:40:@7248.6]
  assign _GEN_1155 = _T_11956 ? 1'h1 : dataKnown_13; // @[StoreQueue.scala 216:40:@7248.6]
  assign _GEN_1156 = initBits_13 ? 1'h0 : _GEN_1151; // @[StoreQueue.scala 204:35:@7215.4]
  assign _GEN_1157 = initBits_13 ? 1'h0 : _GEN_1155; // @[StoreQueue.scala 204:35:@7215.4]
  assign _GEN_1158 = initBits_13 ? addrQ_13 : _GEN_1150; // @[StoreQueue.scala 204:35:@7215.4]
  assign _GEN_1159 = initBits_13 ? dataQ_13 : _GEN_1154; // @[StoreQueue.scala 204:35:@7215.4]
  assign _T_11965 = inputAddrPriorityPorts_0_14 & _T_4420; // @[StoreQueue.scala 209:52:@7261.6]
  assign _T_11966 = _T_11965 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7262.6]
  assign _T_11969 = inputAddrPriorityPorts_1_14 & _T_4420; // @[StoreQueue.scala 209:52:@7264.6]
  assign _T_11970 = _T_11969 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7265.6]
  assign _T_11981 = _T_11966 | _T_11970; // @[StoreQueue.scala 210:30:@7270.6]
  assign _T_11982 = {_T_11970,_T_11966}; // @[OneHot.scala 18:45:@7272.8]
  assign _T_11983 = _T_11982[1]; // @[CircuitMath.scala 30:8:@7273.8]
  assign _GEN_1161 = _T_11983 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7274.8]
  assign _GEN_1162 = _T_11981 ? _GEN_1161 : addrQ_14; // @[StoreQueue.scala 210:40:@7271.6]
  assign _GEN_1163 = _T_11981 ? 1'h1 : addrKnown_14; // @[StoreQueue.scala 210:40:@7271.6]
  assign _T_11988 = inputDataPriorityPorts_0_14 & _T_4490; // @[StoreQueue.scala 215:52:@7278.6]
  assign _T_11989 = _T_11988 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7279.6]
  assign _T_11992 = inputDataPriorityPorts_1_14 & _T_4490; // @[StoreQueue.scala 215:52:@7281.6]
  assign _T_11993 = _T_11992 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7282.6]
  assign _T_12004 = _T_11989 | _T_11993; // @[StoreQueue.scala 216:30:@7287.6]
  assign _T_12005 = {_T_11993,_T_11989}; // @[OneHot.scala 18:45:@7289.8]
  assign _T_12006 = _T_12005[1]; // @[CircuitMath.scala 30:8:@7290.8]
  assign _GEN_1165 = _T_12006 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7291.8]
  assign _GEN_1166 = _T_12004 ? _GEN_1165 : dataQ_14; // @[StoreQueue.scala 216:40:@7288.6]
  assign _GEN_1167 = _T_12004 ? 1'h1 : dataKnown_14; // @[StoreQueue.scala 216:40:@7288.6]
  assign _GEN_1168 = initBits_14 ? 1'h0 : _GEN_1163; // @[StoreQueue.scala 204:35:@7255.4]
  assign _GEN_1169 = initBits_14 ? 1'h0 : _GEN_1167; // @[StoreQueue.scala 204:35:@7255.4]
  assign _GEN_1170 = initBits_14 ? addrQ_14 : _GEN_1162; // @[StoreQueue.scala 204:35:@7255.4]
  assign _GEN_1171 = initBits_14 ? dataQ_14 : _GEN_1166; // @[StoreQueue.scala 204:35:@7255.4]
  assign _T_12013 = inputAddrPriorityPorts_0_15 & _T_4423; // @[StoreQueue.scala 209:52:@7301.6]
  assign _T_12014 = _T_12013 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@7302.6]
  assign _T_12017 = inputAddrPriorityPorts_1_15 & _T_4423; // @[StoreQueue.scala 209:52:@7304.6]
  assign _T_12018 = _T_12017 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@7305.6]
  assign _T_12029 = _T_12014 | _T_12018; // @[StoreQueue.scala 210:30:@7310.6]
  assign _T_12030 = {_T_12018,_T_12014}; // @[OneHot.scala 18:45:@7312.8]
  assign _T_12031 = _T_12030[1]; // @[CircuitMath.scala 30:8:@7313.8]
  assign _GEN_1173 = _T_12031 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@7314.8]
  assign _GEN_1174 = _T_12029 ? _GEN_1173 : addrQ_15; // @[StoreQueue.scala 210:40:@7311.6]
  assign _GEN_1175 = _T_12029 ? 1'h1 : addrKnown_15; // @[StoreQueue.scala 210:40:@7311.6]
  assign _T_12036 = inputDataPriorityPorts_0_15 & _T_4493; // @[StoreQueue.scala 215:52:@7318.6]
  assign _T_12037 = _T_12036 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@7319.6]
  assign _T_12040 = inputDataPriorityPorts_1_15 & _T_4493; // @[StoreQueue.scala 215:52:@7321.6]
  assign _T_12041 = _T_12040 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@7322.6]
  assign _T_12052 = _T_12037 | _T_12041; // @[StoreQueue.scala 216:30:@7327.6]
  assign _T_12053 = {_T_12041,_T_12037}; // @[OneHot.scala 18:45:@7329.8]
  assign _T_12054 = _T_12053[1]; // @[CircuitMath.scala 30:8:@7330.8]
  assign _GEN_1177 = _T_12054 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@7331.8]
  assign _GEN_1178 = _T_12052 ? _GEN_1177 : dataQ_15; // @[StoreQueue.scala 216:40:@7328.6]
  assign _GEN_1179 = _T_12052 ? 1'h1 : dataKnown_15; // @[StoreQueue.scala 216:40:@7328.6]
  assign _GEN_1180 = initBits_15 ? 1'h0 : _GEN_1175; // @[StoreQueue.scala 204:35:@7295.4]
  assign _GEN_1181 = initBits_15 ? 1'h0 : _GEN_1179; // @[StoreQueue.scala 204:35:@7295.4]
  assign _GEN_1182 = initBits_15 ? addrQ_15 : _GEN_1174; // @[StoreQueue.scala 204:35:@7295.4]
  assign _GEN_1183 = initBits_15 ? dataQ_15 : _GEN_1178; // @[StoreQueue.scala 204:35:@7295.4]
  assign _T_12057 = storeRequest & io_memIsReadyForStores; // @[StoreQueue.scala 229:23:@7335.4]
  assign _T_12060 = head + 4'h1; // @[util.scala 10:8:@7337.6]
  assign _GEN_544 = _T_12060 % 5'h10; // @[util.scala 10:14:@7338.6]
  assign _T_12061 = _GEN_544[4:0]; // @[util.scala 10:14:@7338.6]
  assign _GEN_1184 = _T_12057 ? _T_12061 : {{1'd0}, head}; // @[StoreQueue.scala 229:50:@7336.4]
  assign _GEN_1298 = {{3'd0}, io_bbNumStores}; // @[util.scala 10:8:@7342.6]
  assign _T_12063 = tail + _GEN_1298; // @[util.scala 10:8:@7342.6]
  assign _GEN_545 = _T_12063 % 5'h10; // @[util.scala 10:14:@7343.6]
  assign _T_12064 = _GEN_545[4:0]; // @[util.scala 10:14:@7343.6]
  assign _GEN_1185 = io_bbStart ? _T_12064 : {{1'd0}, tail}; // @[StoreQueue.scala 233:20:@7341.4]
  assign _T_12066 = allocatedEntries_0 == 1'h0; // @[StoreQueue.scala 237:84:@7346.4]
  assign _T_12067 = storeCompleted_0 | _T_12066; // @[StoreQueue.scala 237:81:@7347.4]
  assign _T_12069 = allocatedEntries_1 == 1'h0; // @[StoreQueue.scala 237:84:@7348.4]
  assign _T_12070 = storeCompleted_1 | _T_12069; // @[StoreQueue.scala 237:81:@7349.4]
  assign _T_12072 = allocatedEntries_2 == 1'h0; // @[StoreQueue.scala 237:84:@7350.4]
  assign _T_12073 = storeCompleted_2 | _T_12072; // @[StoreQueue.scala 237:81:@7351.4]
  assign _T_12075 = allocatedEntries_3 == 1'h0; // @[StoreQueue.scala 237:84:@7352.4]
  assign _T_12076 = storeCompleted_3 | _T_12075; // @[StoreQueue.scala 237:81:@7353.4]
  assign _T_12078 = allocatedEntries_4 == 1'h0; // @[StoreQueue.scala 237:84:@7354.4]
  assign _T_12079 = storeCompleted_4 | _T_12078; // @[StoreQueue.scala 237:81:@7355.4]
  assign _T_12081 = allocatedEntries_5 == 1'h0; // @[StoreQueue.scala 237:84:@7356.4]
  assign _T_12082 = storeCompleted_5 | _T_12081; // @[StoreQueue.scala 237:81:@7357.4]
  assign _T_12084 = allocatedEntries_6 == 1'h0; // @[StoreQueue.scala 237:84:@7358.4]
  assign _T_12085 = storeCompleted_6 | _T_12084; // @[StoreQueue.scala 237:81:@7359.4]
  assign _T_12087 = allocatedEntries_7 == 1'h0; // @[StoreQueue.scala 237:84:@7360.4]
  assign _T_12088 = storeCompleted_7 | _T_12087; // @[StoreQueue.scala 237:81:@7361.4]
  assign _T_12090 = allocatedEntries_8 == 1'h0; // @[StoreQueue.scala 237:84:@7362.4]
  assign _T_12091 = storeCompleted_8 | _T_12090; // @[StoreQueue.scala 237:81:@7363.4]
  assign _T_12093 = allocatedEntries_9 == 1'h0; // @[StoreQueue.scala 237:84:@7364.4]
  assign _T_12094 = storeCompleted_9 | _T_12093; // @[StoreQueue.scala 237:81:@7365.4]
  assign _T_12096 = allocatedEntries_10 == 1'h0; // @[StoreQueue.scala 237:84:@7366.4]
  assign _T_12097 = storeCompleted_10 | _T_12096; // @[StoreQueue.scala 237:81:@7367.4]
  assign _T_12099 = allocatedEntries_11 == 1'h0; // @[StoreQueue.scala 237:84:@7368.4]
  assign _T_12100 = storeCompleted_11 | _T_12099; // @[StoreQueue.scala 237:81:@7369.4]
  assign _T_12102 = allocatedEntries_12 == 1'h0; // @[StoreQueue.scala 237:84:@7370.4]
  assign _T_12103 = storeCompleted_12 | _T_12102; // @[StoreQueue.scala 237:81:@7371.4]
  assign _T_12105 = allocatedEntries_13 == 1'h0; // @[StoreQueue.scala 237:84:@7372.4]
  assign _T_12106 = storeCompleted_13 | _T_12105; // @[StoreQueue.scala 237:81:@7373.4]
  assign _T_12108 = allocatedEntries_14 == 1'h0; // @[StoreQueue.scala 237:84:@7374.4]
  assign _T_12109 = storeCompleted_14 | _T_12108; // @[StoreQueue.scala 237:81:@7375.4]
  assign _T_12111 = allocatedEntries_15 == 1'h0; // @[StoreQueue.scala 237:84:@7376.4]
  assign _T_12112 = storeCompleted_15 | _T_12111; // @[StoreQueue.scala 237:81:@7377.4]
  assign _T_12137 = _T_12067 & _T_12070; // @[StoreQueue.scala 237:98:@7396.4]
  assign _T_12138 = _T_12137 & _T_12073; // @[StoreQueue.scala 237:98:@7397.4]
  assign _T_12139 = _T_12138 & _T_12076; // @[StoreQueue.scala 237:98:@7398.4]
  assign _T_12140 = _T_12139 & _T_12079; // @[StoreQueue.scala 237:98:@7399.4]
  assign _T_12141 = _T_12140 & _T_12082; // @[StoreQueue.scala 237:98:@7400.4]
  assign _T_12142 = _T_12141 & _T_12085; // @[StoreQueue.scala 237:98:@7401.4]
  assign _T_12143 = _T_12142 & _T_12088; // @[StoreQueue.scala 237:98:@7402.4]
  assign _T_12144 = _T_12143 & _T_12091; // @[StoreQueue.scala 237:98:@7403.4]
  assign _T_12145 = _T_12144 & _T_12094; // @[StoreQueue.scala 237:98:@7404.4]
  assign _T_12146 = _T_12145 & _T_12097; // @[StoreQueue.scala 237:98:@7405.4]
  assign _T_12147 = _T_12146 & _T_12100; // @[StoreQueue.scala 237:98:@7406.4]
  assign _T_12148 = _T_12147 & _T_12103; // @[StoreQueue.scala 237:98:@7407.4]
  assign _T_12149 = _T_12148 & _T_12106; // @[StoreQueue.scala 237:98:@7408.4]
  assign _T_12150 = _T_12149 & _T_12109; // @[StoreQueue.scala 237:98:@7409.4]
  assign _GEN_1187 = 4'h1 == head ? dataQ_1 : dataQ_0; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1188 = 4'h2 == head ? dataQ_2 : _GEN_1187; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1189 = 4'h3 == head ? dataQ_3 : _GEN_1188; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1190 = 4'h4 == head ? dataQ_4 : _GEN_1189; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1191 = 4'h5 == head ? dataQ_5 : _GEN_1190; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1192 = 4'h6 == head ? dataQ_6 : _GEN_1191; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1193 = 4'h7 == head ? dataQ_7 : _GEN_1192; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1194 = 4'h8 == head ? dataQ_8 : _GEN_1193; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1195 = 4'h9 == head ? dataQ_9 : _GEN_1194; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1196 = 4'ha == head ? dataQ_10 : _GEN_1195; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1197 = 4'hb == head ? dataQ_11 : _GEN_1196; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1198 = 4'hc == head ? dataQ_12 : _GEN_1197; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1199 = 4'hd == head ? dataQ_13 : _GEN_1198; // @[StoreQueue.scala 252:21:@7479.4]
  assign _GEN_1200 = 4'he == head ? dataQ_14 : _GEN_1199; // @[StoreQueue.scala 252:21:@7479.4]
  assign io_storeTail = tail; // @[StoreQueue.scala 246:16:@7413.4]
  assign io_storeHead = head; // @[StoreQueue.scala 245:16:@7412.4]
  assign io_storeEmpty = _T_12150 & _T_12112; // @[StoreQueue.scala 237:17:@7411.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[StoreQueue.scala 250:20:@7462.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[StoreQueue.scala 250:20:@7463.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[StoreQueue.scala 250:20:@7464.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[StoreQueue.scala 250:20:@7465.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[StoreQueue.scala 250:20:@7466.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[StoreQueue.scala 250:20:@7467.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[StoreQueue.scala 250:20:@7468.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[StoreQueue.scala 250:20:@7469.4]
  assign io_storeAddrDone_8 = addrKnown_8; // @[StoreQueue.scala 250:20:@7470.4]
  assign io_storeAddrDone_9 = addrKnown_9; // @[StoreQueue.scala 250:20:@7471.4]
  assign io_storeAddrDone_10 = addrKnown_10; // @[StoreQueue.scala 250:20:@7472.4]
  assign io_storeAddrDone_11 = addrKnown_11; // @[StoreQueue.scala 250:20:@7473.4]
  assign io_storeAddrDone_12 = addrKnown_12; // @[StoreQueue.scala 250:20:@7474.4]
  assign io_storeAddrDone_13 = addrKnown_13; // @[StoreQueue.scala 250:20:@7475.4]
  assign io_storeAddrDone_14 = addrKnown_14; // @[StoreQueue.scala 250:20:@7476.4]
  assign io_storeAddrDone_15 = addrKnown_15; // @[StoreQueue.scala 250:20:@7477.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[StoreQueue.scala 249:20:@7446.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[StoreQueue.scala 249:20:@7447.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[StoreQueue.scala 249:20:@7448.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[StoreQueue.scala 249:20:@7449.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[StoreQueue.scala 249:20:@7450.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[StoreQueue.scala 249:20:@7451.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[StoreQueue.scala 249:20:@7452.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[StoreQueue.scala 249:20:@7453.4]
  assign io_storeDataDone_8 = dataKnown_8; // @[StoreQueue.scala 249:20:@7454.4]
  assign io_storeDataDone_9 = dataKnown_9; // @[StoreQueue.scala 249:20:@7455.4]
  assign io_storeDataDone_10 = dataKnown_10; // @[StoreQueue.scala 249:20:@7456.4]
  assign io_storeDataDone_11 = dataKnown_11; // @[StoreQueue.scala 249:20:@7457.4]
  assign io_storeDataDone_12 = dataKnown_12; // @[StoreQueue.scala 249:20:@7458.4]
  assign io_storeDataDone_13 = dataKnown_13; // @[StoreQueue.scala 249:20:@7459.4]
  assign io_storeDataDone_14 = dataKnown_14; // @[StoreQueue.scala 249:20:@7460.4]
  assign io_storeDataDone_15 = dataKnown_15; // @[StoreQueue.scala 249:20:@7461.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[StoreQueue.scala 247:21:@7414.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[StoreQueue.scala 247:21:@7415.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[StoreQueue.scala 247:21:@7416.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[StoreQueue.scala 247:21:@7417.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[StoreQueue.scala 247:21:@7418.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[StoreQueue.scala 247:21:@7419.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[StoreQueue.scala 247:21:@7420.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[StoreQueue.scala 247:21:@7421.4]
  assign io_storeAddrQueue_8 = addrQ_8; // @[StoreQueue.scala 247:21:@7422.4]
  assign io_storeAddrQueue_9 = addrQ_9; // @[StoreQueue.scala 247:21:@7423.4]
  assign io_storeAddrQueue_10 = addrQ_10; // @[StoreQueue.scala 247:21:@7424.4]
  assign io_storeAddrQueue_11 = addrQ_11; // @[StoreQueue.scala 247:21:@7425.4]
  assign io_storeAddrQueue_12 = addrQ_12; // @[StoreQueue.scala 247:21:@7426.4]
  assign io_storeAddrQueue_13 = addrQ_13; // @[StoreQueue.scala 247:21:@7427.4]
  assign io_storeAddrQueue_14 = addrQ_14; // @[StoreQueue.scala 247:21:@7428.4]
  assign io_storeAddrQueue_15 = addrQ_15; // @[StoreQueue.scala 247:21:@7429.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[StoreQueue.scala 248:21:@7430.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[StoreQueue.scala 248:21:@7431.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[StoreQueue.scala 248:21:@7432.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[StoreQueue.scala 248:21:@7433.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[StoreQueue.scala 248:21:@7434.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[StoreQueue.scala 248:21:@7435.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[StoreQueue.scala 248:21:@7436.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[StoreQueue.scala 248:21:@7437.4]
  assign io_storeDataQueue_8 = dataQ_8; // @[StoreQueue.scala 248:21:@7438.4]
  assign io_storeDataQueue_9 = dataQ_9; // @[StoreQueue.scala 248:21:@7439.4]
  assign io_storeDataQueue_10 = dataQ_10; // @[StoreQueue.scala 248:21:@7440.4]
  assign io_storeDataQueue_11 = dataQ_11; // @[StoreQueue.scala 248:21:@7441.4]
  assign io_storeDataQueue_12 = dataQ_12; // @[StoreQueue.scala 248:21:@7442.4]
  assign io_storeDataQueue_13 = dataQ_13; // @[StoreQueue.scala 248:21:@7443.4]
  assign io_storeDataQueue_14 = dataQ_14; // @[StoreQueue.scala 248:21:@7444.4]
  assign io_storeDataQueue_15 = dataQ_15; // @[StoreQueue.scala 248:21:@7445.4]
  assign io_storeAddrToMem = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 253:21:@7480.4]
  assign io_storeDataToMem = 4'hf == head ? dataQ_15 : _GEN_1200; // @[StoreQueue.scala 252:21:@7479.4]
  assign io_storeEnableToMem = _T_3533 & _T_3550; // @[StoreQueue.scala 251:23:@7478.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  storeCompleted_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  storeCompleted_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  storeCompleted_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  storeCompleted_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  storeCompleted_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  storeCompleted_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  storeCompleted_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  storeCompleted_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  checkBits_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  checkBits_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  checkBits_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  checkBits_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  checkBits_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  checkBits_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  checkBits_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  checkBits_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  checkBits_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  checkBits_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  checkBits_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  checkBits_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  checkBits_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  checkBits_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  checkBits_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  checkBits_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  previousLoadHead = _RAND_146[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_1184[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_1185[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1812) begin
          offsetQ_0 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1812) begin
            offsetQ_0 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1812) begin
              offsetQ_0 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1812) begin
                offsetQ_0 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1812) begin
                  offsetQ_0 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1812) begin
                    offsetQ_0 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1812) begin
                      offsetQ_0 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1812) begin
                        offsetQ_0 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1812) begin
                          offsetQ_0 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1812) begin
                            offsetQ_0 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1812) begin
                              offsetQ_0 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1812) begin
                                offsetQ_0 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1812) begin
                                  offsetQ_0 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1812) begin
                                    offsetQ_0 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1812) begin
                                      offsetQ_0 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1830) begin
          offsetQ_1 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1830) begin
            offsetQ_1 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1830) begin
              offsetQ_1 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1830) begin
                offsetQ_1 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1830) begin
                  offsetQ_1 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1830) begin
                    offsetQ_1 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1830) begin
                      offsetQ_1 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1830) begin
                        offsetQ_1 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1830) begin
                          offsetQ_1 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1830) begin
                            offsetQ_1 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1830) begin
                              offsetQ_1 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1830) begin
                                offsetQ_1 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1830) begin
                                  offsetQ_1 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1830) begin
                                    offsetQ_1 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1830) begin
                                      offsetQ_1 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1848) begin
          offsetQ_2 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1848) begin
            offsetQ_2 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1848) begin
              offsetQ_2 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1848) begin
                offsetQ_2 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1848) begin
                  offsetQ_2 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1848) begin
                    offsetQ_2 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1848) begin
                      offsetQ_2 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1848) begin
                        offsetQ_2 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1848) begin
                          offsetQ_2 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1848) begin
                            offsetQ_2 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1848) begin
                              offsetQ_2 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1848) begin
                                offsetQ_2 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1848) begin
                                  offsetQ_2 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1848) begin
                                    offsetQ_2 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1848) begin
                                      offsetQ_2 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1866) begin
          offsetQ_3 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1866) begin
            offsetQ_3 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1866) begin
              offsetQ_3 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1866) begin
                offsetQ_3 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1866) begin
                  offsetQ_3 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1866) begin
                    offsetQ_3 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1866) begin
                      offsetQ_3 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1866) begin
                        offsetQ_3 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1866) begin
                          offsetQ_3 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1866) begin
                            offsetQ_3 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1866) begin
                              offsetQ_3 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1866) begin
                                offsetQ_3 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1866) begin
                                  offsetQ_3 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1866) begin
                                    offsetQ_3 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1866) begin
                                      offsetQ_3 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1884) begin
          offsetQ_4 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1884) begin
            offsetQ_4 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1884) begin
              offsetQ_4 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1884) begin
                offsetQ_4 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1884) begin
                  offsetQ_4 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1884) begin
                    offsetQ_4 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1884) begin
                      offsetQ_4 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1884) begin
                        offsetQ_4 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1884) begin
                          offsetQ_4 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1884) begin
                            offsetQ_4 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1884) begin
                              offsetQ_4 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1884) begin
                                offsetQ_4 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1884) begin
                                  offsetQ_4 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1884) begin
                                    offsetQ_4 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1884) begin
                                      offsetQ_4 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_1902) begin
          offsetQ_5 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1902) begin
            offsetQ_5 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1902) begin
              offsetQ_5 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1902) begin
                offsetQ_5 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1902) begin
                  offsetQ_5 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1902) begin
                    offsetQ_5 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1902) begin
                      offsetQ_5 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1902) begin
                        offsetQ_5 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1902) begin
                          offsetQ_5 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1902) begin
                            offsetQ_5 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1902) begin
                              offsetQ_5 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1902) begin
                                offsetQ_5 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1902) begin
                                  offsetQ_5 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1902) begin
                                    offsetQ_5 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1902) begin
                                      offsetQ_5 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_1920) begin
          offsetQ_6 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1920) begin
            offsetQ_6 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1920) begin
              offsetQ_6 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1920) begin
                offsetQ_6 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1920) begin
                  offsetQ_6 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1920) begin
                    offsetQ_6 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1920) begin
                      offsetQ_6 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1920) begin
                        offsetQ_6 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1920) begin
                          offsetQ_6 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1920) begin
                            offsetQ_6 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1920) begin
                              offsetQ_6 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1920) begin
                                offsetQ_6 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1920) begin
                                  offsetQ_6 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1920) begin
                                    offsetQ_6 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1920) begin
                                      offsetQ_6 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_1938) begin
          offsetQ_7 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1938) begin
            offsetQ_7 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1938) begin
              offsetQ_7 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1938) begin
                offsetQ_7 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1938) begin
                  offsetQ_7 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1938) begin
                    offsetQ_7 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1938) begin
                      offsetQ_7 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1938) begin
                        offsetQ_7 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1938) begin
                          offsetQ_7 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1938) begin
                            offsetQ_7 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1938) begin
                              offsetQ_7 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1938) begin
                                offsetQ_7 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1938) begin
                                  offsetQ_7 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1938) begin
                                    offsetQ_7 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1938) begin
                                      offsetQ_7 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_1956) begin
          offsetQ_8 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1956) begin
            offsetQ_8 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1956) begin
              offsetQ_8 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1956) begin
                offsetQ_8 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1956) begin
                  offsetQ_8 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1956) begin
                    offsetQ_8 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1956) begin
                      offsetQ_8 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1956) begin
                        offsetQ_8 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1956) begin
                          offsetQ_8 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1956) begin
                            offsetQ_8 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1956) begin
                              offsetQ_8 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1956) begin
                                offsetQ_8 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1956) begin
                                  offsetQ_8 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1956) begin
                                    offsetQ_8 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1956) begin
                                      offsetQ_8 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_1974) begin
          offsetQ_9 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1974) begin
            offsetQ_9 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1974) begin
              offsetQ_9 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1974) begin
                offsetQ_9 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1974) begin
                  offsetQ_9 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1974) begin
                    offsetQ_9 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1974) begin
                      offsetQ_9 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1974) begin
                        offsetQ_9 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1974) begin
                          offsetQ_9 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1974) begin
                            offsetQ_9 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1974) begin
                              offsetQ_9 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1974) begin
                                offsetQ_9 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1974) begin
                                  offsetQ_9 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1974) begin
                                    offsetQ_9 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1974) begin
                                      offsetQ_9 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_1992) begin
          offsetQ_10 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1992) begin
            offsetQ_10 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1992) begin
              offsetQ_10 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1992) begin
                offsetQ_10 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1992) begin
                  offsetQ_10 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1992) begin
                    offsetQ_10 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1992) begin
                      offsetQ_10 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1992) begin
                        offsetQ_10 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1992) begin
                          offsetQ_10 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1992) begin
                            offsetQ_10 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1992) begin
                              offsetQ_10 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1992) begin
                                offsetQ_10 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1992) begin
                                  offsetQ_10 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1992) begin
                                    offsetQ_10 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1992) begin
                                      offsetQ_10 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2010) begin
          offsetQ_11 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2010) begin
            offsetQ_11 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2010) begin
              offsetQ_11 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2010) begin
                offsetQ_11 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2010) begin
                  offsetQ_11 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2010) begin
                    offsetQ_11 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2010) begin
                      offsetQ_11 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2010) begin
                        offsetQ_11 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2010) begin
                          offsetQ_11 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2010) begin
                            offsetQ_11 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2010) begin
                              offsetQ_11 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2010) begin
                                offsetQ_11 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2010) begin
                                  offsetQ_11 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2010) begin
                                    offsetQ_11 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2010) begin
                                      offsetQ_11 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2028) begin
          offsetQ_12 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2028) begin
            offsetQ_12 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2028) begin
              offsetQ_12 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2028) begin
                offsetQ_12 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2028) begin
                  offsetQ_12 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2028) begin
                    offsetQ_12 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2028) begin
                      offsetQ_12 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2028) begin
                        offsetQ_12 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2028) begin
                          offsetQ_12 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2028) begin
                            offsetQ_12 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2028) begin
                              offsetQ_12 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2028) begin
                                offsetQ_12 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2028) begin
                                  offsetQ_12 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2028) begin
                                    offsetQ_12 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2028) begin
                                      offsetQ_12 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2046) begin
          offsetQ_13 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2046) begin
            offsetQ_13 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2046) begin
              offsetQ_13 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2046) begin
                offsetQ_13 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2046) begin
                  offsetQ_13 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2046) begin
                    offsetQ_13 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2046) begin
                      offsetQ_13 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2046) begin
                        offsetQ_13 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2046) begin
                          offsetQ_13 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2046) begin
                            offsetQ_13 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2046) begin
                              offsetQ_13 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2046) begin
                                offsetQ_13 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2046) begin
                                  offsetQ_13 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2046) begin
                                    offsetQ_13 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2046) begin
                                      offsetQ_13 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2064) begin
          offsetQ_14 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2064) begin
            offsetQ_14 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2064) begin
              offsetQ_14 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2064) begin
                offsetQ_14 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2064) begin
                  offsetQ_14 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2064) begin
                    offsetQ_14 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2064) begin
                      offsetQ_14 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2064) begin
                        offsetQ_14 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2064) begin
                          offsetQ_14 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2064) begin
                            offsetQ_14 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2064) begin
                              offsetQ_14 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2064) begin
                                offsetQ_14 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2064) begin
                                  offsetQ_14 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2064) begin
                                    offsetQ_14 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2064) begin
                                      offsetQ_14 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2082) begin
          offsetQ_15 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2082) begin
            offsetQ_15 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2082) begin
              offsetQ_15 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2082) begin
                offsetQ_15 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2082) begin
                  offsetQ_15 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2082) begin
                    offsetQ_15 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2082) begin
                      offsetQ_15 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2082) begin
                        offsetQ_15 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2082) begin
                          offsetQ_15 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2082) begin
                            offsetQ_15 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2082) begin
                              offsetQ_15 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2082) begin
                                offsetQ_15 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2082) begin
                                  offsetQ_15 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2082) begin
                                    offsetQ_15 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2082) begin
                                      offsetQ_15 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1812) begin
          portQ_0 <= 1'h0;
        end else begin
          if (4'he == _T_1812) begin
            portQ_0 <= 1'h0;
          end else begin
            if (4'hd == _T_1812) begin
              portQ_0 <= 1'h0;
            end else begin
              if (4'hc == _T_1812) begin
                portQ_0 <= 1'h0;
              end else begin
                if (4'hb == _T_1812) begin
                  portQ_0 <= 1'h0;
                end else begin
                  if (4'ha == _T_1812) begin
                    portQ_0 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1812) begin
                      portQ_0 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1812) begin
                        portQ_0 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1812) begin
                          portQ_0 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1812) begin
                            portQ_0 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1812) begin
                              portQ_0 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1812) begin
                                portQ_0 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1812) begin
                                  portQ_0 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1812) begin
                                    portQ_0 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1812) begin
                                      portQ_0 <= 1'h0;
                                    end else begin
                                      portQ_0 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1830) begin
          portQ_1 <= 1'h0;
        end else begin
          if (4'he == _T_1830) begin
            portQ_1 <= 1'h0;
          end else begin
            if (4'hd == _T_1830) begin
              portQ_1 <= 1'h0;
            end else begin
              if (4'hc == _T_1830) begin
                portQ_1 <= 1'h0;
              end else begin
                if (4'hb == _T_1830) begin
                  portQ_1 <= 1'h0;
                end else begin
                  if (4'ha == _T_1830) begin
                    portQ_1 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1830) begin
                      portQ_1 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1830) begin
                        portQ_1 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1830) begin
                          portQ_1 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1830) begin
                            portQ_1 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1830) begin
                              portQ_1 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1830) begin
                                portQ_1 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1830) begin
                                  portQ_1 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1830) begin
                                    portQ_1 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1830) begin
                                      portQ_1 <= 1'h0;
                                    end else begin
                                      portQ_1 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1848) begin
          portQ_2 <= 1'h0;
        end else begin
          if (4'he == _T_1848) begin
            portQ_2 <= 1'h0;
          end else begin
            if (4'hd == _T_1848) begin
              portQ_2 <= 1'h0;
            end else begin
              if (4'hc == _T_1848) begin
                portQ_2 <= 1'h0;
              end else begin
                if (4'hb == _T_1848) begin
                  portQ_2 <= 1'h0;
                end else begin
                  if (4'ha == _T_1848) begin
                    portQ_2 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1848) begin
                      portQ_2 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1848) begin
                        portQ_2 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1848) begin
                          portQ_2 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1848) begin
                            portQ_2 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1848) begin
                              portQ_2 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1848) begin
                                portQ_2 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1848) begin
                                  portQ_2 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1848) begin
                                    portQ_2 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1848) begin
                                      portQ_2 <= 1'h0;
                                    end else begin
                                      portQ_2 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1866) begin
          portQ_3 <= 1'h0;
        end else begin
          if (4'he == _T_1866) begin
            portQ_3 <= 1'h0;
          end else begin
            if (4'hd == _T_1866) begin
              portQ_3 <= 1'h0;
            end else begin
              if (4'hc == _T_1866) begin
                portQ_3 <= 1'h0;
              end else begin
                if (4'hb == _T_1866) begin
                  portQ_3 <= 1'h0;
                end else begin
                  if (4'ha == _T_1866) begin
                    portQ_3 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1866) begin
                      portQ_3 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1866) begin
                        portQ_3 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1866) begin
                          portQ_3 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1866) begin
                            portQ_3 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1866) begin
                              portQ_3 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1866) begin
                                portQ_3 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1866) begin
                                  portQ_3 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1866) begin
                                    portQ_3 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1866) begin
                                      portQ_3 <= 1'h0;
                                    end else begin
                                      portQ_3 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1884) begin
          portQ_4 <= 1'h0;
        end else begin
          if (4'he == _T_1884) begin
            portQ_4 <= 1'h0;
          end else begin
            if (4'hd == _T_1884) begin
              portQ_4 <= 1'h0;
            end else begin
              if (4'hc == _T_1884) begin
                portQ_4 <= 1'h0;
              end else begin
                if (4'hb == _T_1884) begin
                  portQ_4 <= 1'h0;
                end else begin
                  if (4'ha == _T_1884) begin
                    portQ_4 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1884) begin
                      portQ_4 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1884) begin
                        portQ_4 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1884) begin
                          portQ_4 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1884) begin
                            portQ_4 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1884) begin
                              portQ_4 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1884) begin
                                portQ_4 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1884) begin
                                  portQ_4 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1884) begin
                                    portQ_4 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1884) begin
                                      portQ_4 <= 1'h0;
                                    end else begin
                                      portQ_4 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_1902) begin
          portQ_5 <= 1'h0;
        end else begin
          if (4'he == _T_1902) begin
            portQ_5 <= 1'h0;
          end else begin
            if (4'hd == _T_1902) begin
              portQ_5 <= 1'h0;
            end else begin
              if (4'hc == _T_1902) begin
                portQ_5 <= 1'h0;
              end else begin
                if (4'hb == _T_1902) begin
                  portQ_5 <= 1'h0;
                end else begin
                  if (4'ha == _T_1902) begin
                    portQ_5 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1902) begin
                      portQ_5 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1902) begin
                        portQ_5 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1902) begin
                          portQ_5 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1902) begin
                            portQ_5 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1902) begin
                              portQ_5 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1902) begin
                                portQ_5 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1902) begin
                                  portQ_5 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1902) begin
                                    portQ_5 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1902) begin
                                      portQ_5 <= 1'h0;
                                    end else begin
                                      portQ_5 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_1920) begin
          portQ_6 <= 1'h0;
        end else begin
          if (4'he == _T_1920) begin
            portQ_6 <= 1'h0;
          end else begin
            if (4'hd == _T_1920) begin
              portQ_6 <= 1'h0;
            end else begin
              if (4'hc == _T_1920) begin
                portQ_6 <= 1'h0;
              end else begin
                if (4'hb == _T_1920) begin
                  portQ_6 <= 1'h0;
                end else begin
                  if (4'ha == _T_1920) begin
                    portQ_6 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1920) begin
                      portQ_6 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1920) begin
                        portQ_6 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1920) begin
                          portQ_6 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1920) begin
                            portQ_6 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1920) begin
                              portQ_6 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1920) begin
                                portQ_6 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1920) begin
                                  portQ_6 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1920) begin
                                    portQ_6 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1920) begin
                                      portQ_6 <= 1'h0;
                                    end else begin
                                      portQ_6 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_1938) begin
          portQ_7 <= 1'h0;
        end else begin
          if (4'he == _T_1938) begin
            portQ_7 <= 1'h0;
          end else begin
            if (4'hd == _T_1938) begin
              portQ_7 <= 1'h0;
            end else begin
              if (4'hc == _T_1938) begin
                portQ_7 <= 1'h0;
              end else begin
                if (4'hb == _T_1938) begin
                  portQ_7 <= 1'h0;
                end else begin
                  if (4'ha == _T_1938) begin
                    portQ_7 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1938) begin
                      portQ_7 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1938) begin
                        portQ_7 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1938) begin
                          portQ_7 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1938) begin
                            portQ_7 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1938) begin
                              portQ_7 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1938) begin
                                portQ_7 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1938) begin
                                  portQ_7 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1938) begin
                                    portQ_7 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1938) begin
                                      portQ_7 <= 1'h0;
                                    end else begin
                                      portQ_7 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_1956) begin
          portQ_8 <= 1'h0;
        end else begin
          if (4'he == _T_1956) begin
            portQ_8 <= 1'h0;
          end else begin
            if (4'hd == _T_1956) begin
              portQ_8 <= 1'h0;
            end else begin
              if (4'hc == _T_1956) begin
                portQ_8 <= 1'h0;
              end else begin
                if (4'hb == _T_1956) begin
                  portQ_8 <= 1'h0;
                end else begin
                  if (4'ha == _T_1956) begin
                    portQ_8 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1956) begin
                      portQ_8 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1956) begin
                        portQ_8 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1956) begin
                          portQ_8 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1956) begin
                            portQ_8 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1956) begin
                              portQ_8 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1956) begin
                                portQ_8 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1956) begin
                                  portQ_8 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1956) begin
                                    portQ_8 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1956) begin
                                      portQ_8 <= 1'h0;
                                    end else begin
                                      portQ_8 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_1974) begin
          portQ_9 <= 1'h0;
        end else begin
          if (4'he == _T_1974) begin
            portQ_9 <= 1'h0;
          end else begin
            if (4'hd == _T_1974) begin
              portQ_9 <= 1'h0;
            end else begin
              if (4'hc == _T_1974) begin
                portQ_9 <= 1'h0;
              end else begin
                if (4'hb == _T_1974) begin
                  portQ_9 <= 1'h0;
                end else begin
                  if (4'ha == _T_1974) begin
                    portQ_9 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1974) begin
                      portQ_9 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1974) begin
                        portQ_9 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1974) begin
                          portQ_9 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1974) begin
                            portQ_9 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1974) begin
                              portQ_9 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1974) begin
                                portQ_9 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1974) begin
                                  portQ_9 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1974) begin
                                    portQ_9 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1974) begin
                                      portQ_9 <= 1'h0;
                                    end else begin
                                      portQ_9 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_1992) begin
          portQ_10 <= 1'h0;
        end else begin
          if (4'he == _T_1992) begin
            portQ_10 <= 1'h0;
          end else begin
            if (4'hd == _T_1992) begin
              portQ_10 <= 1'h0;
            end else begin
              if (4'hc == _T_1992) begin
                portQ_10 <= 1'h0;
              end else begin
                if (4'hb == _T_1992) begin
                  portQ_10 <= 1'h0;
                end else begin
                  if (4'ha == _T_1992) begin
                    portQ_10 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_1992) begin
                      portQ_10 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_1992) begin
                        portQ_10 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_1992) begin
                          portQ_10 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_1992) begin
                            portQ_10 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_1992) begin
                              portQ_10 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_1992) begin
                                portQ_10 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_1992) begin
                                  portQ_10 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_1992) begin
                                    portQ_10 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_1992) begin
                                      portQ_10 <= 1'h0;
                                    end else begin
                                      portQ_10 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2010) begin
          portQ_11 <= 1'h0;
        end else begin
          if (4'he == _T_2010) begin
            portQ_11 <= 1'h0;
          end else begin
            if (4'hd == _T_2010) begin
              portQ_11 <= 1'h0;
            end else begin
              if (4'hc == _T_2010) begin
                portQ_11 <= 1'h0;
              end else begin
                if (4'hb == _T_2010) begin
                  portQ_11 <= 1'h0;
                end else begin
                  if (4'ha == _T_2010) begin
                    portQ_11 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2010) begin
                      portQ_11 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2010) begin
                        portQ_11 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2010) begin
                          portQ_11 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2010) begin
                            portQ_11 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2010) begin
                              portQ_11 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2010) begin
                                portQ_11 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2010) begin
                                  portQ_11 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2010) begin
                                    portQ_11 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2010) begin
                                      portQ_11 <= 1'h0;
                                    end else begin
                                      portQ_11 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2028) begin
          portQ_12 <= 1'h0;
        end else begin
          if (4'he == _T_2028) begin
            portQ_12 <= 1'h0;
          end else begin
            if (4'hd == _T_2028) begin
              portQ_12 <= 1'h0;
            end else begin
              if (4'hc == _T_2028) begin
                portQ_12 <= 1'h0;
              end else begin
                if (4'hb == _T_2028) begin
                  portQ_12 <= 1'h0;
                end else begin
                  if (4'ha == _T_2028) begin
                    portQ_12 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2028) begin
                      portQ_12 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2028) begin
                        portQ_12 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2028) begin
                          portQ_12 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2028) begin
                            portQ_12 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2028) begin
                              portQ_12 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2028) begin
                                portQ_12 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2028) begin
                                  portQ_12 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2028) begin
                                    portQ_12 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2028) begin
                                      portQ_12 <= 1'h0;
                                    end else begin
                                      portQ_12 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2046) begin
          portQ_13 <= 1'h0;
        end else begin
          if (4'he == _T_2046) begin
            portQ_13 <= 1'h0;
          end else begin
            if (4'hd == _T_2046) begin
              portQ_13 <= 1'h0;
            end else begin
              if (4'hc == _T_2046) begin
                portQ_13 <= 1'h0;
              end else begin
                if (4'hb == _T_2046) begin
                  portQ_13 <= 1'h0;
                end else begin
                  if (4'ha == _T_2046) begin
                    portQ_13 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2046) begin
                      portQ_13 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2046) begin
                        portQ_13 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2046) begin
                          portQ_13 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2046) begin
                            portQ_13 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2046) begin
                              portQ_13 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2046) begin
                                portQ_13 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2046) begin
                                  portQ_13 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2046) begin
                                    portQ_13 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2046) begin
                                      portQ_13 <= 1'h0;
                                    end else begin
                                      portQ_13 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2064) begin
          portQ_14 <= 1'h0;
        end else begin
          if (4'he == _T_2064) begin
            portQ_14 <= 1'h0;
          end else begin
            if (4'hd == _T_2064) begin
              portQ_14 <= 1'h0;
            end else begin
              if (4'hc == _T_2064) begin
                portQ_14 <= 1'h0;
              end else begin
                if (4'hb == _T_2064) begin
                  portQ_14 <= 1'h0;
                end else begin
                  if (4'ha == _T_2064) begin
                    portQ_14 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2064) begin
                      portQ_14 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2064) begin
                        portQ_14 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2064) begin
                          portQ_14 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2064) begin
                            portQ_14 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2064) begin
                              portQ_14 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2064) begin
                                portQ_14 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2064) begin
                                  portQ_14 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2064) begin
                                    portQ_14 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2064) begin
                                      portQ_14 <= 1'h0;
                                    end else begin
                                      portQ_14 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2082) begin
          portQ_15 <= 1'h0;
        end else begin
          if (4'he == _T_2082) begin
            portQ_15 <= 1'h0;
          end else begin
            if (4'hd == _T_2082) begin
              portQ_15 <= 1'h0;
            end else begin
              if (4'hc == _T_2082) begin
                portQ_15 <= 1'h0;
              end else begin
                if (4'hb == _T_2082) begin
                  portQ_15 <= 1'h0;
                end else begin
                  if (4'ha == _T_2082) begin
                    portQ_15 <= 1'h0;
                  end else begin
                    if (4'h9 == _T_2082) begin
                      portQ_15 <= 1'h0;
                    end else begin
                      if (4'h8 == _T_2082) begin
                        portQ_15 <= 1'h0;
                      end else begin
                        if (4'h7 == _T_2082) begin
                          portQ_15 <= 1'h0;
                        end else begin
                          if (4'h6 == _T_2082) begin
                            portQ_15 <= 1'h0;
                          end else begin
                            if (4'h5 == _T_2082) begin
                              portQ_15 <= 1'h0;
                            end else begin
                              if (4'h4 == _T_2082) begin
                                portQ_15 <= 1'h0;
                              end else begin
                                if (4'h3 == _T_2082) begin
                                  portQ_15 <= 1'h0;
                                end else begin
                                  if (4'h2 == _T_2082) begin
                                    portQ_15 <= 1'h0;
                                  end else begin
                                    if (4'h1 == _T_2082) begin
                                      portQ_15 <= 1'h0;
                                    end else begin
                                      portQ_15 <= io_bbStorePorts_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_11309) begin
          if (_T_11311) begin
            addrQ_0 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_0 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_11357) begin
          if (_T_11359) begin
            addrQ_1 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_1 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_11405) begin
          if (_T_11407) begin
            addrQ_2 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_2 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_11453) begin
          if (_T_11455) begin
            addrQ_3 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_3 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_11501) begin
          if (_T_11503) begin
            addrQ_4 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_4 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_11549) begin
          if (_T_11551) begin
            addrQ_5 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_5 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_11597) begin
          if (_T_11599) begin
            addrQ_6 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_6 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_11645) begin
          if (_T_11647) begin
            addrQ_7 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_7 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_11693) begin
          if (_T_11695) begin
            addrQ_8 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_8 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_11741) begin
          if (_T_11743) begin
            addrQ_9 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_9 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_11789) begin
          if (_T_11791) begin
            addrQ_10 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_10 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_11837) begin
          if (_T_11839) begin
            addrQ_11 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_11 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_11885) begin
          if (_T_11887) begin
            addrQ_12 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_12 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_11933) begin
          if (_T_11935) begin
            addrQ_13 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_13 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_11981) begin
          if (_T_11983) begin
            addrQ_14 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_14 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_12029) begin
          if (_T_12031) begin
            addrQ_15 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_15 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_11332) begin
          if (_T_11334) begin
            dataQ_0 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_0 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_11380) begin
          if (_T_11382) begin
            dataQ_1 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_1 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_11428) begin
          if (_T_11430) begin
            dataQ_2 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_2 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_11476) begin
          if (_T_11478) begin
            dataQ_3 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_3 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_11524) begin
          if (_T_11526) begin
            dataQ_4 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_4 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_11572) begin
          if (_T_11574) begin
            dataQ_5 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_5 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_11620) begin
          if (_T_11622) begin
            dataQ_6 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_6 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_11668) begin
          if (_T_11670) begin
            dataQ_7 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_7 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_11716) begin
          if (_T_11718) begin
            dataQ_8 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_8 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_11764) begin
          if (_T_11766) begin
            dataQ_9 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_9 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_11812) begin
          if (_T_11814) begin
            dataQ_10 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_10 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_11860) begin
          if (_T_11862) begin
            dataQ_11 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_11 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_11908) begin
          if (_T_11910) begin
            dataQ_12 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_12 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_11956) begin
          if (_T_11958) begin
            dataQ_13 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_13 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_12004) begin
          if (_T_12006) begin
            dataQ_14 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_14 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_12052) begin
          if (_T_12054) begin
            dataQ_15 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_15 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_11309) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_11357) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_11405) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_11453) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_11501) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_11549) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_11597) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_11645) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_11693) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_11741) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_11789) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_11837) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_11885) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_11933) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_11981) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_12029) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_11332) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_11380) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_11428) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_11476) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_11524) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_11572) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_11620) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_11668) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_11716) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_11764) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_11812) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_11860) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_11908) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_11956) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_12004) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_12052) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1766;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1767;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1768;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1769;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1770;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1771;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1772;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1773;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1774;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1775;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1776;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1777;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1778;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1779;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1780;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1781;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_3555) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_3561) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_3567) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_3573) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_3579) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_3585) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_3591) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_3597) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        storeCompleted_8 <= 1'h0;
      end else begin
        if (_T_3603) begin
          storeCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        storeCompleted_9 <= 1'h0;
      end else begin
        if (_T_3609) begin
          storeCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        storeCompleted_10 <= 1'h0;
      end else begin
        if (_T_3615) begin
          storeCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        storeCompleted_11 <= 1'h0;
      end else begin
        if (_T_3621) begin
          storeCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        storeCompleted_12 <= 1'h0;
      end else begin
        if (_T_3627) begin
          storeCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        storeCompleted_13 <= 1'h0;
      end else begin
        if (_T_3633) begin
          storeCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        storeCompleted_14 <= 1'h0;
      end else begin
        if (_T_3639) begin
          storeCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        storeCompleted_15 <= 1'h0;
      end else begin
        if (_T_3645) begin
          storeCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2109;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2113) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2121) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2139;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2143) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2151) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2169;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2173) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2181) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2199;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2203) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2211) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2229;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2233) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2241) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2259;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2263) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2271) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2289;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2293) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2301) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2319;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2323) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2331) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2349;
      end else begin
        if (io_loadEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2353) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2361) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2379;
      end else begin
        if (io_loadEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2383) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2391) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2409;
      end else begin
        if (io_loadEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2413) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2421) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2439;
      end else begin
        if (io_loadEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2443) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2451) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2469;
      end else begin
        if (io_loadEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2473) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2481) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2499;
      end else begin
        if (io_loadEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2503) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2511) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2529;
      end else begin
        if (io_loadEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2533) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2541) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2559;
      end else begin
        if (io_loadEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2563) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2571) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_E( // @[:@7482.2]
  input         clock, // @[:@7483.4]
  input         reset, // @[:@7484.4]
  input         io_bbStart, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_0, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_1, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_2, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_3, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_4, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_5, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_6, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_7, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_8, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_9, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_10, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_11, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_12, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_13, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_14, // @[:@7485.4]
  input  [3:0]  io_bbLoadOffsets_15, // @[:@7485.4]
  input         io_bbNumLoads, // @[:@7485.4]
  output [3:0]  io_loadTail, // @[:@7485.4]
  output [3:0]  io_loadHead, // @[:@7485.4]
  output        io_loadEmpty, // @[:@7485.4]
  input  [3:0]  io_storeTail, // @[:@7485.4]
  input  [3:0]  io_storeHead, // @[:@7485.4]
  input         io_storeEmpty, // @[:@7485.4]
  input         io_storeAddrDone_0, // @[:@7485.4]
  input         io_storeAddrDone_1, // @[:@7485.4]
  input         io_storeAddrDone_2, // @[:@7485.4]
  input         io_storeAddrDone_3, // @[:@7485.4]
  input         io_storeAddrDone_4, // @[:@7485.4]
  input         io_storeAddrDone_5, // @[:@7485.4]
  input         io_storeAddrDone_6, // @[:@7485.4]
  input         io_storeAddrDone_7, // @[:@7485.4]
  input         io_storeAddrDone_8, // @[:@7485.4]
  input         io_storeAddrDone_9, // @[:@7485.4]
  input         io_storeAddrDone_10, // @[:@7485.4]
  input         io_storeAddrDone_11, // @[:@7485.4]
  input         io_storeAddrDone_12, // @[:@7485.4]
  input         io_storeAddrDone_13, // @[:@7485.4]
  input         io_storeAddrDone_14, // @[:@7485.4]
  input         io_storeAddrDone_15, // @[:@7485.4]
  input         io_storeDataDone_0, // @[:@7485.4]
  input         io_storeDataDone_1, // @[:@7485.4]
  input         io_storeDataDone_2, // @[:@7485.4]
  input         io_storeDataDone_3, // @[:@7485.4]
  input         io_storeDataDone_4, // @[:@7485.4]
  input         io_storeDataDone_5, // @[:@7485.4]
  input         io_storeDataDone_6, // @[:@7485.4]
  input         io_storeDataDone_7, // @[:@7485.4]
  input         io_storeDataDone_8, // @[:@7485.4]
  input         io_storeDataDone_9, // @[:@7485.4]
  input         io_storeDataDone_10, // @[:@7485.4]
  input         io_storeDataDone_11, // @[:@7485.4]
  input         io_storeDataDone_12, // @[:@7485.4]
  input         io_storeDataDone_13, // @[:@7485.4]
  input         io_storeDataDone_14, // @[:@7485.4]
  input         io_storeDataDone_15, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_0, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_1, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_2, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_3, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_4, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_5, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_6, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_7, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_8, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_9, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_10, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_11, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_12, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_13, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_14, // @[:@7485.4]
  input  [31:0] io_storeAddrQueue_15, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_0, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_1, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_2, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_3, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_4, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_5, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_6, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_7, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_8, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_9, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_10, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_11, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_12, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_13, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_14, // @[:@7485.4]
  input  [31:0] io_storeDataQueue_15, // @[:@7485.4]
  output        io_loadAddrDone_0, // @[:@7485.4]
  output        io_loadAddrDone_1, // @[:@7485.4]
  output        io_loadAddrDone_2, // @[:@7485.4]
  output        io_loadAddrDone_3, // @[:@7485.4]
  output        io_loadAddrDone_4, // @[:@7485.4]
  output        io_loadAddrDone_5, // @[:@7485.4]
  output        io_loadAddrDone_6, // @[:@7485.4]
  output        io_loadAddrDone_7, // @[:@7485.4]
  output        io_loadAddrDone_8, // @[:@7485.4]
  output        io_loadAddrDone_9, // @[:@7485.4]
  output        io_loadAddrDone_10, // @[:@7485.4]
  output        io_loadAddrDone_11, // @[:@7485.4]
  output        io_loadAddrDone_12, // @[:@7485.4]
  output        io_loadAddrDone_13, // @[:@7485.4]
  output        io_loadAddrDone_14, // @[:@7485.4]
  output        io_loadAddrDone_15, // @[:@7485.4]
  output        io_loadDataDone_0, // @[:@7485.4]
  output        io_loadDataDone_1, // @[:@7485.4]
  output        io_loadDataDone_2, // @[:@7485.4]
  output        io_loadDataDone_3, // @[:@7485.4]
  output        io_loadDataDone_4, // @[:@7485.4]
  output        io_loadDataDone_5, // @[:@7485.4]
  output        io_loadDataDone_6, // @[:@7485.4]
  output        io_loadDataDone_7, // @[:@7485.4]
  output        io_loadDataDone_8, // @[:@7485.4]
  output        io_loadDataDone_9, // @[:@7485.4]
  output        io_loadDataDone_10, // @[:@7485.4]
  output        io_loadDataDone_11, // @[:@7485.4]
  output        io_loadDataDone_12, // @[:@7485.4]
  output        io_loadDataDone_13, // @[:@7485.4]
  output        io_loadDataDone_14, // @[:@7485.4]
  output        io_loadDataDone_15, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_0, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_1, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_2, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_3, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_4, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_5, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_6, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_7, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_8, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_9, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_10, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_11, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_12, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_13, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_14, // @[:@7485.4]
  output [31:0] io_loadAddrQueue_15, // @[:@7485.4]
  input         io_loadAddrEnable_0, // @[:@7485.4]
  input  [31:0] io_addrFromLoadPorts_0, // @[:@7485.4]
  input         io_loadPorts_0_ready, // @[:@7485.4]
  output        io_loadPorts_0_valid, // @[:@7485.4]
  output [31:0] io_loadPorts_0_bits, // @[:@7485.4]
  input  [31:0] io_loadDataFromMem, // @[:@7485.4]
  output [31:0] io_loadAddrToMem, // @[:@7485.4]
  output        io_loadEnableToMem, // @[:@7485.4]
  input         io_memIsReadyForLoads // @[:@7485.4]
);
  reg [3:0] head; // @[LoadQueue.scala 50:21:@7487.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[LoadQueue.scala 51:21:@7488.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[LoadQueue.scala 53:24:@7506.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[LoadQueue.scala 54:22:@7524.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[LoadQueue.scala 55:22:@7542.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[LoadQueue.scala 56:22:@7560.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[LoadQueue.scala 57:26:@7578.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[LoadQueue.scala 58:26:@7596.4]
  reg [31:0] _RAND_97;
  reg  loadCompleted_0; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_98;
  reg  loadCompleted_1; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_99;
  reg  loadCompleted_2; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_100;
  reg  loadCompleted_3; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_101;
  reg  loadCompleted_4; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_102;
  reg  loadCompleted_5; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_103;
  reg  loadCompleted_6; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_104;
  reg  loadCompleted_7; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_105;
  reg  loadCompleted_8; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_106;
  reg  loadCompleted_9; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_107;
  reg  loadCompleted_10; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_108;
  reg  loadCompleted_11; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_109;
  reg  loadCompleted_12; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_110;
  reg  loadCompleted_13; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_111;
  reg  loadCompleted_14; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_112;
  reg  loadCompleted_15; // @[LoadQueue.scala 59:30:@7614.4]
  reg [31:0] _RAND_113;
  reg  allocatedEntries_0; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_114;
  reg  allocatedEntries_1; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_115;
  reg  allocatedEntries_2; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_116;
  reg  allocatedEntries_3; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_117;
  reg  allocatedEntries_4; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_118;
  reg  allocatedEntries_5; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_119;
  reg  allocatedEntries_6; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_120;
  reg  allocatedEntries_7; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_121;
  reg  allocatedEntries_8; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_122;
  reg  allocatedEntries_9; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_123;
  reg  allocatedEntries_10; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_124;
  reg  allocatedEntries_11; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_125;
  reg  allocatedEntries_12; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_126;
  reg  allocatedEntries_13; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_127;
  reg  allocatedEntries_14; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_128;
  reg  allocatedEntries_15; // @[LoadQueue.scala 60:33:@7632.4]
  reg [31:0] _RAND_129;
  reg  bypassInitiated_0; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_130;
  reg  bypassInitiated_1; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_131;
  reg  bypassInitiated_2; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_132;
  reg  bypassInitiated_3; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_133;
  reg  bypassInitiated_4; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_134;
  reg  bypassInitiated_5; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_135;
  reg  bypassInitiated_6; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_136;
  reg  bypassInitiated_7; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_137;
  reg  bypassInitiated_8; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_138;
  reg  bypassInitiated_9; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_139;
  reg  bypassInitiated_10; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_140;
  reg  bypassInitiated_11; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_141;
  reg  bypassInitiated_12; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_142;
  reg  bypassInitiated_13; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_143;
  reg  bypassInitiated_14; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_144;
  reg  bypassInitiated_15; // @[LoadQueue.scala 61:32:@7650.4]
  reg [31:0] _RAND_145;
  reg  checkBits_0; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_146;
  reg  checkBits_1; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_147;
  reg  checkBits_2; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_148;
  reg  checkBits_3; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_149;
  reg  checkBits_4; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_150;
  reg  checkBits_5; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_151;
  reg  checkBits_6; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_152;
  reg  checkBits_7; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_153;
  reg  checkBits_8; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_154;
  reg  checkBits_9; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_155;
  reg  checkBits_10; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_156;
  reg  checkBits_11; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_157;
  reg  checkBits_12; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_158;
  reg  checkBits_13; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_159;
  reg  checkBits_14; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_160;
  reg  checkBits_15; // @[LoadQueue.scala 62:26:@7668.4]
  reg [31:0] _RAND_161;
  wire [5:0] _GEN_2262; // @[util.scala 14:20:@7670.4]
  wire [6:0] _T_1716; // @[util.scala 14:20:@7670.4]
  wire [6:0] _T_1717; // @[util.scala 14:20:@7671.4]
  wire [5:0] _T_1718; // @[util.scala 14:20:@7672.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@7673.4]
  wire [4:0] _T_1719; // @[util.scala 14:25:@7673.4]
  wire [4:0] _GEN_2263; // @[LoadQueue.scala 71:46:@7674.4]
  wire  _T_1720; // @[LoadQueue.scala 71:46:@7674.4]
  wire  initBits_0; // @[LoadQueue.scala 71:63:@7675.4]
  wire [6:0] _T_1725; // @[util.scala 14:20:@7677.4]
  wire [6:0] _T_1726; // @[util.scala 14:20:@7678.4]
  wire [5:0] _T_1727; // @[util.scala 14:20:@7679.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@7680.4]
  wire [4:0] _T_1728; // @[util.scala 14:25:@7680.4]
  wire  _T_1729; // @[LoadQueue.scala 71:46:@7681.4]
  wire  initBits_1; // @[LoadQueue.scala 71:63:@7682.4]
  wire [6:0] _T_1734; // @[util.scala 14:20:@7684.4]
  wire [6:0] _T_1735; // @[util.scala 14:20:@7685.4]
  wire [5:0] _T_1736; // @[util.scala 14:20:@7686.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@7687.4]
  wire [4:0] _T_1737; // @[util.scala 14:25:@7687.4]
  wire  _T_1738; // @[LoadQueue.scala 71:46:@7688.4]
  wire  initBits_2; // @[LoadQueue.scala 71:63:@7689.4]
  wire [6:0] _T_1743; // @[util.scala 14:20:@7691.4]
  wire [6:0] _T_1744; // @[util.scala 14:20:@7692.4]
  wire [5:0] _T_1745; // @[util.scala 14:20:@7693.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@7694.4]
  wire [4:0] _T_1746; // @[util.scala 14:25:@7694.4]
  wire  _T_1747; // @[LoadQueue.scala 71:46:@7695.4]
  wire  initBits_3; // @[LoadQueue.scala 71:63:@7696.4]
  wire [6:0] _T_1752; // @[util.scala 14:20:@7698.4]
  wire [6:0] _T_1753; // @[util.scala 14:20:@7699.4]
  wire [5:0] _T_1754; // @[util.scala 14:20:@7700.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@7701.4]
  wire [4:0] _T_1755; // @[util.scala 14:25:@7701.4]
  wire  _T_1756; // @[LoadQueue.scala 71:46:@7702.4]
  wire  initBits_4; // @[LoadQueue.scala 71:63:@7703.4]
  wire [6:0] _T_1761; // @[util.scala 14:20:@7705.4]
  wire [6:0] _T_1762; // @[util.scala 14:20:@7706.4]
  wire [5:0] _T_1763; // @[util.scala 14:20:@7707.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@7708.4]
  wire [4:0] _T_1764; // @[util.scala 14:25:@7708.4]
  wire  _T_1765; // @[LoadQueue.scala 71:46:@7709.4]
  wire  initBits_5; // @[LoadQueue.scala 71:63:@7710.4]
  wire [6:0] _T_1770; // @[util.scala 14:20:@7712.4]
  wire [6:0] _T_1771; // @[util.scala 14:20:@7713.4]
  wire [5:0] _T_1772; // @[util.scala 14:20:@7714.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@7715.4]
  wire [4:0] _T_1773; // @[util.scala 14:25:@7715.4]
  wire  _T_1774; // @[LoadQueue.scala 71:46:@7716.4]
  wire  initBits_6; // @[LoadQueue.scala 71:63:@7717.4]
  wire [6:0] _T_1779; // @[util.scala 14:20:@7719.4]
  wire [6:0] _T_1780; // @[util.scala 14:20:@7720.4]
  wire [5:0] _T_1781; // @[util.scala 14:20:@7721.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@7722.4]
  wire [4:0] _T_1782; // @[util.scala 14:25:@7722.4]
  wire  _T_1783; // @[LoadQueue.scala 71:46:@7723.4]
  wire  initBits_7; // @[LoadQueue.scala 71:63:@7724.4]
  wire [6:0] _T_1788; // @[util.scala 14:20:@7726.4]
  wire [6:0] _T_1789; // @[util.scala 14:20:@7727.4]
  wire [5:0] _T_1790; // @[util.scala 14:20:@7728.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@7729.4]
  wire [4:0] _T_1791; // @[util.scala 14:25:@7729.4]
  wire  _T_1792; // @[LoadQueue.scala 71:46:@7730.4]
  wire  initBits_8; // @[LoadQueue.scala 71:63:@7731.4]
  wire [6:0] _T_1797; // @[util.scala 14:20:@7733.4]
  wire [6:0] _T_1798; // @[util.scala 14:20:@7734.4]
  wire [5:0] _T_1799; // @[util.scala 14:20:@7735.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@7736.4]
  wire [4:0] _T_1800; // @[util.scala 14:25:@7736.4]
  wire  _T_1801; // @[LoadQueue.scala 71:46:@7737.4]
  wire  initBits_9; // @[LoadQueue.scala 71:63:@7738.4]
  wire [6:0] _T_1806; // @[util.scala 14:20:@7740.4]
  wire [6:0] _T_1807; // @[util.scala 14:20:@7741.4]
  wire [5:0] _T_1808; // @[util.scala 14:20:@7742.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@7743.4]
  wire [4:0] _T_1809; // @[util.scala 14:25:@7743.4]
  wire  _T_1810; // @[LoadQueue.scala 71:46:@7744.4]
  wire  initBits_10; // @[LoadQueue.scala 71:63:@7745.4]
  wire [6:0] _T_1815; // @[util.scala 14:20:@7747.4]
  wire [6:0] _T_1816; // @[util.scala 14:20:@7748.4]
  wire [5:0] _T_1817; // @[util.scala 14:20:@7749.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@7750.4]
  wire [4:0] _T_1818; // @[util.scala 14:25:@7750.4]
  wire  _T_1819; // @[LoadQueue.scala 71:46:@7751.4]
  wire  initBits_11; // @[LoadQueue.scala 71:63:@7752.4]
  wire [6:0] _T_1824; // @[util.scala 14:20:@7754.4]
  wire [6:0] _T_1825; // @[util.scala 14:20:@7755.4]
  wire [5:0] _T_1826; // @[util.scala 14:20:@7756.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@7757.4]
  wire [4:0] _T_1827; // @[util.scala 14:25:@7757.4]
  wire  _T_1828; // @[LoadQueue.scala 71:46:@7758.4]
  wire  initBits_12; // @[LoadQueue.scala 71:63:@7759.4]
  wire [6:0] _T_1833; // @[util.scala 14:20:@7761.4]
  wire [6:0] _T_1834; // @[util.scala 14:20:@7762.4]
  wire [5:0] _T_1835; // @[util.scala 14:20:@7763.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@7764.4]
  wire [4:0] _T_1836; // @[util.scala 14:25:@7764.4]
  wire  _T_1837; // @[LoadQueue.scala 71:46:@7765.4]
  wire  initBits_13; // @[LoadQueue.scala 71:63:@7766.4]
  wire [6:0] _T_1842; // @[util.scala 14:20:@7768.4]
  wire [6:0] _T_1843; // @[util.scala 14:20:@7769.4]
  wire [5:0] _T_1844; // @[util.scala 14:20:@7770.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@7771.4]
  wire [4:0] _T_1845; // @[util.scala 14:25:@7771.4]
  wire  _T_1846; // @[LoadQueue.scala 71:46:@7772.4]
  wire  initBits_14; // @[LoadQueue.scala 71:63:@7773.4]
  wire [6:0] _T_1851; // @[util.scala 14:20:@7775.4]
  wire [6:0] _T_1852; // @[util.scala 14:20:@7776.4]
  wire [5:0] _T_1853; // @[util.scala 14:20:@7777.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@7778.4]
  wire [4:0] _T_1854; // @[util.scala 14:25:@7778.4]
  wire  _T_1855; // @[LoadQueue.scala 71:46:@7779.4]
  wire  initBits_15; // @[LoadQueue.scala 71:63:@7780.4]
  wire  _T_1878; // @[LoadQueue.scala 73:78:@7798.4]
  wire  _T_1879; // @[LoadQueue.scala 73:78:@7799.4]
  wire  _T_1880; // @[LoadQueue.scala 73:78:@7800.4]
  wire  _T_1881; // @[LoadQueue.scala 73:78:@7801.4]
  wire  _T_1882; // @[LoadQueue.scala 73:78:@7802.4]
  wire  _T_1883; // @[LoadQueue.scala 73:78:@7803.4]
  wire  _T_1884; // @[LoadQueue.scala 73:78:@7804.4]
  wire  _T_1885; // @[LoadQueue.scala 73:78:@7805.4]
  wire  _T_1886; // @[LoadQueue.scala 73:78:@7806.4]
  wire  _T_1887; // @[LoadQueue.scala 73:78:@7807.4]
  wire  _T_1888; // @[LoadQueue.scala 73:78:@7808.4]
  wire  _T_1889; // @[LoadQueue.scala 73:78:@7809.4]
  wire  _T_1890; // @[LoadQueue.scala 73:78:@7810.4]
  wire  _T_1891; // @[LoadQueue.scala 73:78:@7811.4]
  wire  _T_1892; // @[LoadQueue.scala 73:78:@7812.4]
  wire  _T_1893; // @[LoadQueue.scala 73:78:@7813.4]
  wire [3:0] _T_1924; // @[:@7853.6]
  wire [3:0] _GEN_1; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_2; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_3; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_4; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_5; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_6; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_7; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_8; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_9; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_10; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_11; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_12; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_13; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_14; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_15; // @[LoadQueue.scala 77:20:@7854.6]
  wire [3:0] _GEN_32; // @[LoadQueue.scala 76:25:@7847.4]
  wire  _GEN_33; // @[LoadQueue.scala 76:25:@7847.4]
  wire [3:0] _T_1942; // @[:@7869.6]
  wire [3:0] _GEN_35; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_36; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_37; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_38; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_39; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_40; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_41; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_42; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_43; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_44; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_45; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_46; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_47; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_48; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_49; // @[LoadQueue.scala 77:20:@7870.6]
  wire [3:0] _GEN_66; // @[LoadQueue.scala 76:25:@7863.4]
  wire  _GEN_67; // @[LoadQueue.scala 76:25:@7863.4]
  wire [3:0] _T_1960; // @[:@7885.6]
  wire [3:0] _GEN_69; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_70; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_71; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_72; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_73; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_74; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_75; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_76; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_77; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_78; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_79; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_80; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_81; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_82; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_83; // @[LoadQueue.scala 77:20:@7886.6]
  wire [3:0] _GEN_100; // @[LoadQueue.scala 76:25:@7879.4]
  wire  _GEN_101; // @[LoadQueue.scala 76:25:@7879.4]
  wire [3:0] _T_1978; // @[:@7901.6]
  wire [3:0] _GEN_103; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_104; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_105; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_106; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_107; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_108; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_109; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_110; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_111; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_112; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_113; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_114; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_115; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_116; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_117; // @[LoadQueue.scala 77:20:@7902.6]
  wire [3:0] _GEN_134; // @[LoadQueue.scala 76:25:@7895.4]
  wire  _GEN_135; // @[LoadQueue.scala 76:25:@7895.4]
  wire [3:0] _T_1996; // @[:@7917.6]
  wire [3:0] _GEN_137; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_138; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_139; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_140; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_141; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_142; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_143; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_144; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_145; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_146; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_147; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_148; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_149; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_150; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_151; // @[LoadQueue.scala 77:20:@7918.6]
  wire [3:0] _GEN_168; // @[LoadQueue.scala 76:25:@7911.4]
  wire  _GEN_169; // @[LoadQueue.scala 76:25:@7911.4]
  wire [3:0] _T_2014; // @[:@7933.6]
  wire [3:0] _GEN_171; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_172; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_173; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_174; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_175; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_176; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_177; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_178; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_179; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_180; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_181; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_182; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_183; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_184; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_185; // @[LoadQueue.scala 77:20:@7934.6]
  wire [3:0] _GEN_202; // @[LoadQueue.scala 76:25:@7927.4]
  wire  _GEN_203; // @[LoadQueue.scala 76:25:@7927.4]
  wire [3:0] _T_2032; // @[:@7949.6]
  wire [3:0] _GEN_205; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_206; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_207; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_208; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_209; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_210; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_211; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_212; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_213; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_214; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_215; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_216; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_217; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_218; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_219; // @[LoadQueue.scala 77:20:@7950.6]
  wire [3:0] _GEN_236; // @[LoadQueue.scala 76:25:@7943.4]
  wire  _GEN_237; // @[LoadQueue.scala 76:25:@7943.4]
  wire [3:0] _T_2050; // @[:@7965.6]
  wire [3:0] _GEN_239; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_240; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_241; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_242; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_243; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_244; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_245; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_246; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_247; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_248; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_249; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_250; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_251; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_252; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_253; // @[LoadQueue.scala 77:20:@7966.6]
  wire [3:0] _GEN_270; // @[LoadQueue.scala 76:25:@7959.4]
  wire  _GEN_271; // @[LoadQueue.scala 76:25:@7959.4]
  wire [3:0] _T_2068; // @[:@7981.6]
  wire [3:0] _GEN_273; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_274; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_275; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_276; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_277; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_278; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_279; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_280; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_281; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_282; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_283; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_284; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_285; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_286; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_287; // @[LoadQueue.scala 77:20:@7982.6]
  wire [3:0] _GEN_304; // @[LoadQueue.scala 76:25:@7975.4]
  wire  _GEN_305; // @[LoadQueue.scala 76:25:@7975.4]
  wire [3:0] _T_2086; // @[:@7997.6]
  wire [3:0] _GEN_307; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_308; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_309; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_310; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_311; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_312; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_313; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_314; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_315; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_316; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_317; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_318; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_319; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_320; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_321; // @[LoadQueue.scala 77:20:@7998.6]
  wire [3:0] _GEN_338; // @[LoadQueue.scala 76:25:@7991.4]
  wire  _GEN_339; // @[LoadQueue.scala 76:25:@7991.4]
  wire [3:0] _T_2104; // @[:@8013.6]
  wire [3:0] _GEN_341; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_342; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_343; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_344; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_345; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_346; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_347; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_348; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_349; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_350; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_351; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_352; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_353; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_354; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_355; // @[LoadQueue.scala 77:20:@8014.6]
  wire [3:0] _GEN_372; // @[LoadQueue.scala 76:25:@8007.4]
  wire  _GEN_373; // @[LoadQueue.scala 76:25:@8007.4]
  wire [3:0] _T_2122; // @[:@8029.6]
  wire [3:0] _GEN_375; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_376; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_377; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_378; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_379; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_380; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_381; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_382; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_383; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_384; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_385; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_386; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_387; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_388; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_389; // @[LoadQueue.scala 77:20:@8030.6]
  wire [3:0] _GEN_406; // @[LoadQueue.scala 76:25:@8023.4]
  wire  _GEN_407; // @[LoadQueue.scala 76:25:@8023.4]
  wire [3:0] _T_2140; // @[:@8045.6]
  wire [3:0] _GEN_409; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_410; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_411; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_412; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_413; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_414; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_415; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_416; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_417; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_418; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_419; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_420; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_421; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_422; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_423; // @[LoadQueue.scala 77:20:@8046.6]
  wire [3:0] _GEN_440; // @[LoadQueue.scala 76:25:@8039.4]
  wire  _GEN_441; // @[LoadQueue.scala 76:25:@8039.4]
  wire [3:0] _T_2158; // @[:@8061.6]
  wire [3:0] _GEN_443; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_444; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_445; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_446; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_447; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_448; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_449; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_450; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_451; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_452; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_453; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_454; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_455; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_456; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_457; // @[LoadQueue.scala 77:20:@8062.6]
  wire [3:0] _GEN_474; // @[LoadQueue.scala 76:25:@8055.4]
  wire  _GEN_475; // @[LoadQueue.scala 76:25:@8055.4]
  wire [3:0] _T_2176; // @[:@8077.6]
  wire [3:0] _GEN_477; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_478; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_479; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_480; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_481; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_482; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_483; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_484; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_485; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_486; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_487; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_488; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_489; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_490; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_491; // @[LoadQueue.scala 77:20:@8078.6]
  wire [3:0] _GEN_508; // @[LoadQueue.scala 76:25:@8071.4]
  wire  _GEN_509; // @[LoadQueue.scala 76:25:@8071.4]
  wire [3:0] _T_2194; // @[:@8093.6]
  wire [3:0] _GEN_511; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_512; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_513; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_514; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_515; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_516; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_517; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_518; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_519; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_520; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_521; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_522; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_523; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_524; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_525; // @[LoadQueue.scala 77:20:@8094.6]
  wire [3:0] _GEN_542; // @[LoadQueue.scala 76:25:@8087.4]
  wire  _GEN_543; // @[LoadQueue.scala 76:25:@8087.4]
  reg [3:0] previousStoreHead; // @[LoadQueue.scala 93:34:@8103.4]
  reg [31:0] _RAND_162;
  wire [4:0] _T_2216; // @[util.scala 10:8:@8112.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@8113.6]
  wire [4:0] _T_2217; // @[util.scala 10:14:@8113.6]
  wire [4:0] _GEN_2327; // @[LoadQueue.scala 97:56:@8114.6]
  wire  _T_2218; // @[LoadQueue.scala 97:56:@8114.6]
  wire  _T_2219; // @[LoadQueue.scala 96:50:@8115.6]
  wire  _T_2221; // @[LoadQueue.scala 96:34:@8116.6]
  wire  _T_2223; // @[LoadQueue.scala 101:36:@8124.8]
  wire  _T_2224; // @[LoadQueue.scala 101:86:@8125.8]
  wire  _T_2225; // @[LoadQueue.scala 101:61:@8126.8]
  wire  _T_2227; // @[LoadQueue.scala 103:36:@8131.10]
  wire  _T_2228; // @[LoadQueue.scala 103:69:@8132.10]
  wire  _T_2229; // @[LoadQueue.scala 104:31:@8133.10]
  wire  _T_2230; // @[LoadQueue.scala 103:94:@8134.10]
  wire  _T_2232; // @[LoadQueue.scala 103:54:@8135.10]
  wire  _T_2233; // @[LoadQueue.scala 103:51:@8136.10]
  wire  _GEN_560; // @[LoadQueue.scala 104:53:@8137.10]
  wire  _GEN_561; // @[LoadQueue.scala 101:102:@8127.8]
  wire  _GEN_562; // @[LoadQueue.scala 99:27:@8120.6]
  wire  _GEN_563; // @[LoadQueue.scala 95:34:@8105.4]
  wire [4:0] _T_2246; // @[util.scala 10:8:@8148.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@8149.6]
  wire [4:0] _T_2247; // @[util.scala 10:14:@8149.6]
  wire  _T_2248; // @[LoadQueue.scala 97:56:@8150.6]
  wire  _T_2249; // @[LoadQueue.scala 96:50:@8151.6]
  wire  _T_2251; // @[LoadQueue.scala 96:34:@8152.6]
  wire  _T_2253; // @[LoadQueue.scala 101:36:@8160.8]
  wire  _T_2254; // @[LoadQueue.scala 101:86:@8161.8]
  wire  _T_2255; // @[LoadQueue.scala 101:61:@8162.8]
  wire  _T_2258; // @[LoadQueue.scala 103:69:@8168.10]
  wire  _T_2259; // @[LoadQueue.scala 104:31:@8169.10]
  wire  _T_2260; // @[LoadQueue.scala 103:94:@8170.10]
  wire  _T_2262; // @[LoadQueue.scala 103:54:@8171.10]
  wire  _T_2263; // @[LoadQueue.scala 103:51:@8172.10]
  wire  _GEN_580; // @[LoadQueue.scala 104:53:@8173.10]
  wire  _GEN_581; // @[LoadQueue.scala 101:102:@8163.8]
  wire  _GEN_582; // @[LoadQueue.scala 99:27:@8156.6]
  wire  _GEN_583; // @[LoadQueue.scala 95:34:@8141.4]
  wire [4:0] _T_2276; // @[util.scala 10:8:@8184.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@8185.6]
  wire [4:0] _T_2277; // @[util.scala 10:14:@8185.6]
  wire  _T_2278; // @[LoadQueue.scala 97:56:@8186.6]
  wire  _T_2279; // @[LoadQueue.scala 96:50:@8187.6]
  wire  _T_2281; // @[LoadQueue.scala 96:34:@8188.6]
  wire  _T_2283; // @[LoadQueue.scala 101:36:@8196.8]
  wire  _T_2284; // @[LoadQueue.scala 101:86:@8197.8]
  wire  _T_2285; // @[LoadQueue.scala 101:61:@8198.8]
  wire  _T_2288; // @[LoadQueue.scala 103:69:@8204.10]
  wire  _T_2289; // @[LoadQueue.scala 104:31:@8205.10]
  wire  _T_2290; // @[LoadQueue.scala 103:94:@8206.10]
  wire  _T_2292; // @[LoadQueue.scala 103:54:@8207.10]
  wire  _T_2293; // @[LoadQueue.scala 103:51:@8208.10]
  wire  _GEN_600; // @[LoadQueue.scala 104:53:@8209.10]
  wire  _GEN_601; // @[LoadQueue.scala 101:102:@8199.8]
  wire  _GEN_602; // @[LoadQueue.scala 99:27:@8192.6]
  wire  _GEN_603; // @[LoadQueue.scala 95:34:@8177.4]
  wire [4:0] _T_2306; // @[util.scala 10:8:@8220.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@8221.6]
  wire [4:0] _T_2307; // @[util.scala 10:14:@8221.6]
  wire  _T_2308; // @[LoadQueue.scala 97:56:@8222.6]
  wire  _T_2309; // @[LoadQueue.scala 96:50:@8223.6]
  wire  _T_2311; // @[LoadQueue.scala 96:34:@8224.6]
  wire  _T_2313; // @[LoadQueue.scala 101:36:@8232.8]
  wire  _T_2314; // @[LoadQueue.scala 101:86:@8233.8]
  wire  _T_2315; // @[LoadQueue.scala 101:61:@8234.8]
  wire  _T_2318; // @[LoadQueue.scala 103:69:@8240.10]
  wire  _T_2319; // @[LoadQueue.scala 104:31:@8241.10]
  wire  _T_2320; // @[LoadQueue.scala 103:94:@8242.10]
  wire  _T_2322; // @[LoadQueue.scala 103:54:@8243.10]
  wire  _T_2323; // @[LoadQueue.scala 103:51:@8244.10]
  wire  _GEN_620; // @[LoadQueue.scala 104:53:@8245.10]
  wire  _GEN_621; // @[LoadQueue.scala 101:102:@8235.8]
  wire  _GEN_622; // @[LoadQueue.scala 99:27:@8228.6]
  wire  _GEN_623; // @[LoadQueue.scala 95:34:@8213.4]
  wire [4:0] _T_2336; // @[util.scala 10:8:@8256.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@8257.6]
  wire [4:0] _T_2337; // @[util.scala 10:14:@8257.6]
  wire  _T_2338; // @[LoadQueue.scala 97:56:@8258.6]
  wire  _T_2339; // @[LoadQueue.scala 96:50:@8259.6]
  wire  _T_2341; // @[LoadQueue.scala 96:34:@8260.6]
  wire  _T_2343; // @[LoadQueue.scala 101:36:@8268.8]
  wire  _T_2344; // @[LoadQueue.scala 101:86:@8269.8]
  wire  _T_2345; // @[LoadQueue.scala 101:61:@8270.8]
  wire  _T_2348; // @[LoadQueue.scala 103:69:@8276.10]
  wire  _T_2349; // @[LoadQueue.scala 104:31:@8277.10]
  wire  _T_2350; // @[LoadQueue.scala 103:94:@8278.10]
  wire  _T_2352; // @[LoadQueue.scala 103:54:@8279.10]
  wire  _T_2353; // @[LoadQueue.scala 103:51:@8280.10]
  wire  _GEN_640; // @[LoadQueue.scala 104:53:@8281.10]
  wire  _GEN_641; // @[LoadQueue.scala 101:102:@8271.8]
  wire  _GEN_642; // @[LoadQueue.scala 99:27:@8264.6]
  wire  _GEN_643; // @[LoadQueue.scala 95:34:@8249.4]
  wire [4:0] _T_2366; // @[util.scala 10:8:@8292.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@8293.6]
  wire [4:0] _T_2367; // @[util.scala 10:14:@8293.6]
  wire  _T_2368; // @[LoadQueue.scala 97:56:@8294.6]
  wire  _T_2369; // @[LoadQueue.scala 96:50:@8295.6]
  wire  _T_2371; // @[LoadQueue.scala 96:34:@8296.6]
  wire  _T_2373; // @[LoadQueue.scala 101:36:@8304.8]
  wire  _T_2374; // @[LoadQueue.scala 101:86:@8305.8]
  wire  _T_2375; // @[LoadQueue.scala 101:61:@8306.8]
  wire  _T_2378; // @[LoadQueue.scala 103:69:@8312.10]
  wire  _T_2379; // @[LoadQueue.scala 104:31:@8313.10]
  wire  _T_2380; // @[LoadQueue.scala 103:94:@8314.10]
  wire  _T_2382; // @[LoadQueue.scala 103:54:@8315.10]
  wire  _T_2383; // @[LoadQueue.scala 103:51:@8316.10]
  wire  _GEN_660; // @[LoadQueue.scala 104:53:@8317.10]
  wire  _GEN_661; // @[LoadQueue.scala 101:102:@8307.8]
  wire  _GEN_662; // @[LoadQueue.scala 99:27:@8300.6]
  wire  _GEN_663; // @[LoadQueue.scala 95:34:@8285.4]
  wire [4:0] _T_2396; // @[util.scala 10:8:@8328.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@8329.6]
  wire [4:0] _T_2397; // @[util.scala 10:14:@8329.6]
  wire  _T_2398; // @[LoadQueue.scala 97:56:@8330.6]
  wire  _T_2399; // @[LoadQueue.scala 96:50:@8331.6]
  wire  _T_2401; // @[LoadQueue.scala 96:34:@8332.6]
  wire  _T_2403; // @[LoadQueue.scala 101:36:@8340.8]
  wire  _T_2404; // @[LoadQueue.scala 101:86:@8341.8]
  wire  _T_2405; // @[LoadQueue.scala 101:61:@8342.8]
  wire  _T_2408; // @[LoadQueue.scala 103:69:@8348.10]
  wire  _T_2409; // @[LoadQueue.scala 104:31:@8349.10]
  wire  _T_2410; // @[LoadQueue.scala 103:94:@8350.10]
  wire  _T_2412; // @[LoadQueue.scala 103:54:@8351.10]
  wire  _T_2413; // @[LoadQueue.scala 103:51:@8352.10]
  wire  _GEN_680; // @[LoadQueue.scala 104:53:@8353.10]
  wire  _GEN_681; // @[LoadQueue.scala 101:102:@8343.8]
  wire  _GEN_682; // @[LoadQueue.scala 99:27:@8336.6]
  wire  _GEN_683; // @[LoadQueue.scala 95:34:@8321.4]
  wire [4:0] _T_2426; // @[util.scala 10:8:@8364.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@8365.6]
  wire [4:0] _T_2427; // @[util.scala 10:14:@8365.6]
  wire  _T_2428; // @[LoadQueue.scala 97:56:@8366.6]
  wire  _T_2429; // @[LoadQueue.scala 96:50:@8367.6]
  wire  _T_2431; // @[LoadQueue.scala 96:34:@8368.6]
  wire  _T_2433; // @[LoadQueue.scala 101:36:@8376.8]
  wire  _T_2434; // @[LoadQueue.scala 101:86:@8377.8]
  wire  _T_2435; // @[LoadQueue.scala 101:61:@8378.8]
  wire  _T_2438; // @[LoadQueue.scala 103:69:@8384.10]
  wire  _T_2439; // @[LoadQueue.scala 104:31:@8385.10]
  wire  _T_2440; // @[LoadQueue.scala 103:94:@8386.10]
  wire  _T_2442; // @[LoadQueue.scala 103:54:@8387.10]
  wire  _T_2443; // @[LoadQueue.scala 103:51:@8388.10]
  wire  _GEN_700; // @[LoadQueue.scala 104:53:@8389.10]
  wire  _GEN_701; // @[LoadQueue.scala 101:102:@8379.8]
  wire  _GEN_702; // @[LoadQueue.scala 99:27:@8372.6]
  wire  _GEN_703; // @[LoadQueue.scala 95:34:@8357.4]
  wire [4:0] _T_2456; // @[util.scala 10:8:@8400.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@8401.6]
  wire [4:0] _T_2457; // @[util.scala 10:14:@8401.6]
  wire  _T_2458; // @[LoadQueue.scala 97:56:@8402.6]
  wire  _T_2459; // @[LoadQueue.scala 96:50:@8403.6]
  wire  _T_2461; // @[LoadQueue.scala 96:34:@8404.6]
  wire  _T_2463; // @[LoadQueue.scala 101:36:@8412.8]
  wire  _T_2464; // @[LoadQueue.scala 101:86:@8413.8]
  wire  _T_2465; // @[LoadQueue.scala 101:61:@8414.8]
  wire  _T_2468; // @[LoadQueue.scala 103:69:@8420.10]
  wire  _T_2469; // @[LoadQueue.scala 104:31:@8421.10]
  wire  _T_2470; // @[LoadQueue.scala 103:94:@8422.10]
  wire  _T_2472; // @[LoadQueue.scala 103:54:@8423.10]
  wire  _T_2473; // @[LoadQueue.scala 103:51:@8424.10]
  wire  _GEN_720; // @[LoadQueue.scala 104:53:@8425.10]
  wire  _GEN_721; // @[LoadQueue.scala 101:102:@8415.8]
  wire  _GEN_722; // @[LoadQueue.scala 99:27:@8408.6]
  wire  _GEN_723; // @[LoadQueue.scala 95:34:@8393.4]
  wire [4:0] _T_2486; // @[util.scala 10:8:@8436.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@8437.6]
  wire [4:0] _T_2487; // @[util.scala 10:14:@8437.6]
  wire  _T_2488; // @[LoadQueue.scala 97:56:@8438.6]
  wire  _T_2489; // @[LoadQueue.scala 96:50:@8439.6]
  wire  _T_2491; // @[LoadQueue.scala 96:34:@8440.6]
  wire  _T_2493; // @[LoadQueue.scala 101:36:@8448.8]
  wire  _T_2494; // @[LoadQueue.scala 101:86:@8449.8]
  wire  _T_2495; // @[LoadQueue.scala 101:61:@8450.8]
  wire  _T_2498; // @[LoadQueue.scala 103:69:@8456.10]
  wire  _T_2499; // @[LoadQueue.scala 104:31:@8457.10]
  wire  _T_2500; // @[LoadQueue.scala 103:94:@8458.10]
  wire  _T_2502; // @[LoadQueue.scala 103:54:@8459.10]
  wire  _T_2503; // @[LoadQueue.scala 103:51:@8460.10]
  wire  _GEN_740; // @[LoadQueue.scala 104:53:@8461.10]
  wire  _GEN_741; // @[LoadQueue.scala 101:102:@8451.8]
  wire  _GEN_742; // @[LoadQueue.scala 99:27:@8444.6]
  wire  _GEN_743; // @[LoadQueue.scala 95:34:@8429.4]
  wire [4:0] _T_2516; // @[util.scala 10:8:@8472.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@8473.6]
  wire [4:0] _T_2517; // @[util.scala 10:14:@8473.6]
  wire  _T_2518; // @[LoadQueue.scala 97:56:@8474.6]
  wire  _T_2519; // @[LoadQueue.scala 96:50:@8475.6]
  wire  _T_2521; // @[LoadQueue.scala 96:34:@8476.6]
  wire  _T_2523; // @[LoadQueue.scala 101:36:@8484.8]
  wire  _T_2524; // @[LoadQueue.scala 101:86:@8485.8]
  wire  _T_2525; // @[LoadQueue.scala 101:61:@8486.8]
  wire  _T_2528; // @[LoadQueue.scala 103:69:@8492.10]
  wire  _T_2529; // @[LoadQueue.scala 104:31:@8493.10]
  wire  _T_2530; // @[LoadQueue.scala 103:94:@8494.10]
  wire  _T_2532; // @[LoadQueue.scala 103:54:@8495.10]
  wire  _T_2533; // @[LoadQueue.scala 103:51:@8496.10]
  wire  _GEN_760; // @[LoadQueue.scala 104:53:@8497.10]
  wire  _GEN_761; // @[LoadQueue.scala 101:102:@8487.8]
  wire  _GEN_762; // @[LoadQueue.scala 99:27:@8480.6]
  wire  _GEN_763; // @[LoadQueue.scala 95:34:@8465.4]
  wire [4:0] _T_2546; // @[util.scala 10:8:@8508.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@8509.6]
  wire [4:0] _T_2547; // @[util.scala 10:14:@8509.6]
  wire  _T_2548; // @[LoadQueue.scala 97:56:@8510.6]
  wire  _T_2549; // @[LoadQueue.scala 96:50:@8511.6]
  wire  _T_2551; // @[LoadQueue.scala 96:34:@8512.6]
  wire  _T_2553; // @[LoadQueue.scala 101:36:@8520.8]
  wire  _T_2554; // @[LoadQueue.scala 101:86:@8521.8]
  wire  _T_2555; // @[LoadQueue.scala 101:61:@8522.8]
  wire  _T_2558; // @[LoadQueue.scala 103:69:@8528.10]
  wire  _T_2559; // @[LoadQueue.scala 104:31:@8529.10]
  wire  _T_2560; // @[LoadQueue.scala 103:94:@8530.10]
  wire  _T_2562; // @[LoadQueue.scala 103:54:@8531.10]
  wire  _T_2563; // @[LoadQueue.scala 103:51:@8532.10]
  wire  _GEN_780; // @[LoadQueue.scala 104:53:@8533.10]
  wire  _GEN_781; // @[LoadQueue.scala 101:102:@8523.8]
  wire  _GEN_782; // @[LoadQueue.scala 99:27:@8516.6]
  wire  _GEN_783; // @[LoadQueue.scala 95:34:@8501.4]
  wire [4:0] _T_2576; // @[util.scala 10:8:@8544.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@8545.6]
  wire [4:0] _T_2577; // @[util.scala 10:14:@8545.6]
  wire  _T_2578; // @[LoadQueue.scala 97:56:@8546.6]
  wire  _T_2579; // @[LoadQueue.scala 96:50:@8547.6]
  wire  _T_2581; // @[LoadQueue.scala 96:34:@8548.6]
  wire  _T_2583; // @[LoadQueue.scala 101:36:@8556.8]
  wire  _T_2584; // @[LoadQueue.scala 101:86:@8557.8]
  wire  _T_2585; // @[LoadQueue.scala 101:61:@8558.8]
  wire  _T_2588; // @[LoadQueue.scala 103:69:@8564.10]
  wire  _T_2589; // @[LoadQueue.scala 104:31:@8565.10]
  wire  _T_2590; // @[LoadQueue.scala 103:94:@8566.10]
  wire  _T_2592; // @[LoadQueue.scala 103:54:@8567.10]
  wire  _T_2593; // @[LoadQueue.scala 103:51:@8568.10]
  wire  _GEN_800; // @[LoadQueue.scala 104:53:@8569.10]
  wire  _GEN_801; // @[LoadQueue.scala 101:102:@8559.8]
  wire  _GEN_802; // @[LoadQueue.scala 99:27:@8552.6]
  wire  _GEN_803; // @[LoadQueue.scala 95:34:@8537.4]
  wire [4:0] _T_2606; // @[util.scala 10:8:@8580.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@8581.6]
  wire [4:0] _T_2607; // @[util.scala 10:14:@8581.6]
  wire  _T_2608; // @[LoadQueue.scala 97:56:@8582.6]
  wire  _T_2609; // @[LoadQueue.scala 96:50:@8583.6]
  wire  _T_2611; // @[LoadQueue.scala 96:34:@8584.6]
  wire  _T_2613; // @[LoadQueue.scala 101:36:@8592.8]
  wire  _T_2614; // @[LoadQueue.scala 101:86:@8593.8]
  wire  _T_2615; // @[LoadQueue.scala 101:61:@8594.8]
  wire  _T_2618; // @[LoadQueue.scala 103:69:@8600.10]
  wire  _T_2619; // @[LoadQueue.scala 104:31:@8601.10]
  wire  _T_2620; // @[LoadQueue.scala 103:94:@8602.10]
  wire  _T_2622; // @[LoadQueue.scala 103:54:@8603.10]
  wire  _T_2623; // @[LoadQueue.scala 103:51:@8604.10]
  wire  _GEN_820; // @[LoadQueue.scala 104:53:@8605.10]
  wire  _GEN_821; // @[LoadQueue.scala 101:102:@8595.8]
  wire  _GEN_822; // @[LoadQueue.scala 99:27:@8588.6]
  wire  _GEN_823; // @[LoadQueue.scala 95:34:@8573.4]
  wire [4:0] _T_2636; // @[util.scala 10:8:@8616.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@8617.6]
  wire [4:0] _T_2637; // @[util.scala 10:14:@8617.6]
  wire  _T_2638; // @[LoadQueue.scala 97:56:@8618.6]
  wire  _T_2639; // @[LoadQueue.scala 96:50:@8619.6]
  wire  _T_2641; // @[LoadQueue.scala 96:34:@8620.6]
  wire  _T_2643; // @[LoadQueue.scala 101:36:@8628.8]
  wire  _T_2644; // @[LoadQueue.scala 101:86:@8629.8]
  wire  _T_2645; // @[LoadQueue.scala 101:61:@8630.8]
  wire  _T_2648; // @[LoadQueue.scala 103:69:@8636.10]
  wire  _T_2649; // @[LoadQueue.scala 104:31:@8637.10]
  wire  _T_2650; // @[LoadQueue.scala 103:94:@8638.10]
  wire  _T_2652; // @[LoadQueue.scala 103:54:@8639.10]
  wire  _T_2653; // @[LoadQueue.scala 103:51:@8640.10]
  wire  _GEN_840; // @[LoadQueue.scala 104:53:@8641.10]
  wire  _GEN_841; // @[LoadQueue.scala 101:102:@8631.8]
  wire  _GEN_842; // @[LoadQueue.scala 99:27:@8624.6]
  wire  _GEN_843; // @[LoadQueue.scala 95:34:@8609.4]
  wire [4:0] _T_2666; // @[util.scala 10:8:@8652.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@8653.6]
  wire [4:0] _T_2667; // @[util.scala 10:14:@8653.6]
  wire  _T_2668; // @[LoadQueue.scala 97:56:@8654.6]
  wire  _T_2669; // @[LoadQueue.scala 96:50:@8655.6]
  wire  _T_2671; // @[LoadQueue.scala 96:34:@8656.6]
  wire  _T_2673; // @[LoadQueue.scala 101:36:@8664.8]
  wire  _T_2674; // @[LoadQueue.scala 101:86:@8665.8]
  wire  _T_2675; // @[LoadQueue.scala 101:61:@8666.8]
  wire  _T_2678; // @[LoadQueue.scala 103:69:@8672.10]
  wire  _T_2679; // @[LoadQueue.scala 104:31:@8673.10]
  wire  _T_2680; // @[LoadQueue.scala 103:94:@8674.10]
  wire  _T_2682; // @[LoadQueue.scala 103:54:@8675.10]
  wire  _T_2683; // @[LoadQueue.scala 103:51:@8676.10]
  wire  _GEN_860; // @[LoadQueue.scala 104:53:@8677.10]
  wire  _GEN_861; // @[LoadQueue.scala 101:102:@8667.8]
  wire  _GEN_862; // @[LoadQueue.scala 99:27:@8660.6]
  wire  _GEN_863; // @[LoadQueue.scala 95:34:@8645.4]
  wire [15:0] _T_2687; // @[OneHot.scala 52:12:@8682.4]
  wire  _T_2689; // @[util.scala 60:60:@8684.4]
  wire  _T_2690; // @[util.scala 60:60:@8685.4]
  wire  _T_2691; // @[util.scala 60:60:@8686.4]
  wire  _T_2692; // @[util.scala 60:60:@8687.4]
  wire  _T_2693; // @[util.scala 60:60:@8688.4]
  wire  _T_2694; // @[util.scala 60:60:@8689.4]
  wire  _T_2695; // @[util.scala 60:60:@8690.4]
  wire  _T_2696; // @[util.scala 60:60:@8691.4]
  wire  _T_2697; // @[util.scala 60:60:@8692.4]
  wire  _T_2698; // @[util.scala 60:60:@8693.4]
  wire  _T_2699; // @[util.scala 60:60:@8694.4]
  wire  _T_2700; // @[util.scala 60:60:@8695.4]
  wire  _T_2701; // @[util.scala 60:60:@8696.4]
  wire  _T_2702; // @[util.scala 60:60:@8697.4]
  wire  _T_2703; // @[util.scala 60:60:@8698.4]
  wire  _T_2704; // @[util.scala 60:60:@8699.4]
  wire [255:0] _T_4835; // @[Mux.scala 19:72:@10223.4]
  wire [255:0] _T_4842; // @[Mux.scala 19:72:@10230.4]
  wire [511:0] _T_4843; // @[Mux.scala 19:72:@10231.4]
  wire [511:0] _T_4845; // @[Mux.scala 19:72:@10232.4]
  wire [255:0] _T_4852; // @[Mux.scala 19:72:@10239.4]
  wire [255:0] _T_4859; // @[Mux.scala 19:72:@10246.4]
  wire [511:0] _T_4860; // @[Mux.scala 19:72:@10247.4]
  wire [511:0] _T_4862; // @[Mux.scala 19:72:@10248.4]
  wire [255:0] _T_4869; // @[Mux.scala 19:72:@10255.4]
  wire [255:0] _T_4876; // @[Mux.scala 19:72:@10262.4]
  wire [511:0] _T_4877; // @[Mux.scala 19:72:@10263.4]
  wire [511:0] _T_4879; // @[Mux.scala 19:72:@10264.4]
  wire [255:0] _T_4886; // @[Mux.scala 19:72:@10271.4]
  wire [255:0] _T_4893; // @[Mux.scala 19:72:@10278.4]
  wire [511:0] _T_4894; // @[Mux.scala 19:72:@10279.4]
  wire [511:0] _T_4896; // @[Mux.scala 19:72:@10280.4]
  wire [255:0] _T_4903; // @[Mux.scala 19:72:@10287.4]
  wire [255:0] _T_4910; // @[Mux.scala 19:72:@10294.4]
  wire [511:0] _T_4911; // @[Mux.scala 19:72:@10295.4]
  wire [511:0] _T_4913; // @[Mux.scala 19:72:@10296.4]
  wire [255:0] _T_4920; // @[Mux.scala 19:72:@10303.4]
  wire [255:0] _T_4927; // @[Mux.scala 19:72:@10310.4]
  wire [511:0] _T_4928; // @[Mux.scala 19:72:@10311.4]
  wire [511:0] _T_4930; // @[Mux.scala 19:72:@10312.4]
  wire [255:0] _T_4937; // @[Mux.scala 19:72:@10319.4]
  wire [255:0] _T_4944; // @[Mux.scala 19:72:@10326.4]
  wire [511:0] _T_4945; // @[Mux.scala 19:72:@10327.4]
  wire [511:0] _T_4947; // @[Mux.scala 19:72:@10328.4]
  wire [255:0] _T_4954; // @[Mux.scala 19:72:@10335.4]
  wire [255:0] _T_4961; // @[Mux.scala 19:72:@10342.4]
  wire [511:0] _T_4962; // @[Mux.scala 19:72:@10343.4]
  wire [511:0] _T_4964; // @[Mux.scala 19:72:@10344.4]
  wire [511:0] _T_4979; // @[Mux.scala 19:72:@10359.4]
  wire [511:0] _T_4981; // @[Mux.scala 19:72:@10360.4]
  wire [511:0] _T_4996; // @[Mux.scala 19:72:@10375.4]
  wire [511:0] _T_4998; // @[Mux.scala 19:72:@10376.4]
  wire [511:0] _T_5013; // @[Mux.scala 19:72:@10391.4]
  wire [511:0] _T_5015; // @[Mux.scala 19:72:@10392.4]
  wire [511:0] _T_5030; // @[Mux.scala 19:72:@10407.4]
  wire [511:0] _T_5032; // @[Mux.scala 19:72:@10408.4]
  wire [511:0] _T_5047; // @[Mux.scala 19:72:@10423.4]
  wire [511:0] _T_5049; // @[Mux.scala 19:72:@10424.4]
  wire [511:0] _T_5064; // @[Mux.scala 19:72:@10439.4]
  wire [511:0] _T_5066; // @[Mux.scala 19:72:@10440.4]
  wire [511:0] _T_5081; // @[Mux.scala 19:72:@10455.4]
  wire [511:0] _T_5083; // @[Mux.scala 19:72:@10456.4]
  wire [511:0] _T_5098; // @[Mux.scala 19:72:@10471.4]
  wire [511:0] _T_5100; // @[Mux.scala 19:72:@10472.4]
  wire [511:0] _T_5101; // @[Mux.scala 19:72:@10473.4]
  wire [511:0] _T_5102; // @[Mux.scala 19:72:@10474.4]
  wire [511:0] _T_5103; // @[Mux.scala 19:72:@10475.4]
  wire [511:0] _T_5104; // @[Mux.scala 19:72:@10476.4]
  wire [511:0] _T_5105; // @[Mux.scala 19:72:@10477.4]
  wire [511:0] _T_5106; // @[Mux.scala 19:72:@10478.4]
  wire [511:0] _T_5107; // @[Mux.scala 19:72:@10479.4]
  wire [511:0] _T_5108; // @[Mux.scala 19:72:@10480.4]
  wire [511:0] _T_5109; // @[Mux.scala 19:72:@10481.4]
  wire [511:0] _T_5110; // @[Mux.scala 19:72:@10482.4]
  wire [511:0] _T_5111; // @[Mux.scala 19:72:@10483.4]
  wire [511:0] _T_5112; // @[Mux.scala 19:72:@10484.4]
  wire [511:0] _T_5113; // @[Mux.scala 19:72:@10485.4]
  wire [511:0] _T_5114; // @[Mux.scala 19:72:@10486.4]
  wire [511:0] _T_5115; // @[Mux.scala 19:72:@10487.4]
  wire [7:0] _T_5692; // @[Mux.scala 19:72:@10837.4]
  wire [7:0] _T_5699; // @[Mux.scala 19:72:@10844.4]
  wire [15:0] _T_5700; // @[Mux.scala 19:72:@10845.4]
  wire [15:0] _T_5702; // @[Mux.scala 19:72:@10846.4]
  wire [7:0] _T_5709; // @[Mux.scala 19:72:@10853.4]
  wire [7:0] _T_5716; // @[Mux.scala 19:72:@10860.4]
  wire [15:0] _T_5717; // @[Mux.scala 19:72:@10861.4]
  wire [15:0] _T_5719; // @[Mux.scala 19:72:@10862.4]
  wire [7:0] _T_5726; // @[Mux.scala 19:72:@10869.4]
  wire [7:0] _T_5733; // @[Mux.scala 19:72:@10876.4]
  wire [15:0] _T_5734; // @[Mux.scala 19:72:@10877.4]
  wire [15:0] _T_5736; // @[Mux.scala 19:72:@10878.4]
  wire [7:0] _T_5743; // @[Mux.scala 19:72:@10885.4]
  wire [7:0] _T_5750; // @[Mux.scala 19:72:@10892.4]
  wire [15:0] _T_5751; // @[Mux.scala 19:72:@10893.4]
  wire [15:0] _T_5753; // @[Mux.scala 19:72:@10894.4]
  wire [7:0] _T_5760; // @[Mux.scala 19:72:@10901.4]
  wire [7:0] _T_5767; // @[Mux.scala 19:72:@10908.4]
  wire [15:0] _T_5768; // @[Mux.scala 19:72:@10909.4]
  wire [15:0] _T_5770; // @[Mux.scala 19:72:@10910.4]
  wire [7:0] _T_5777; // @[Mux.scala 19:72:@10917.4]
  wire [7:0] _T_5784; // @[Mux.scala 19:72:@10924.4]
  wire [15:0] _T_5785; // @[Mux.scala 19:72:@10925.4]
  wire [15:0] _T_5787; // @[Mux.scala 19:72:@10926.4]
  wire [7:0] _T_5794; // @[Mux.scala 19:72:@10933.4]
  wire [7:0] _T_5801; // @[Mux.scala 19:72:@10940.4]
  wire [15:0] _T_5802; // @[Mux.scala 19:72:@10941.4]
  wire [15:0] _T_5804; // @[Mux.scala 19:72:@10942.4]
  wire [7:0] _T_5811; // @[Mux.scala 19:72:@10949.4]
  wire [7:0] _T_5818; // @[Mux.scala 19:72:@10956.4]
  wire [15:0] _T_5819; // @[Mux.scala 19:72:@10957.4]
  wire [15:0] _T_5821; // @[Mux.scala 19:72:@10958.4]
  wire [15:0] _T_5836; // @[Mux.scala 19:72:@10973.4]
  wire [15:0] _T_5838; // @[Mux.scala 19:72:@10974.4]
  wire [15:0] _T_5853; // @[Mux.scala 19:72:@10989.4]
  wire [15:0] _T_5855; // @[Mux.scala 19:72:@10990.4]
  wire [15:0] _T_5870; // @[Mux.scala 19:72:@11005.4]
  wire [15:0] _T_5872; // @[Mux.scala 19:72:@11006.4]
  wire [15:0] _T_5887; // @[Mux.scala 19:72:@11021.4]
  wire [15:0] _T_5889; // @[Mux.scala 19:72:@11022.4]
  wire [15:0] _T_5904; // @[Mux.scala 19:72:@11037.4]
  wire [15:0] _T_5906; // @[Mux.scala 19:72:@11038.4]
  wire [15:0] _T_5921; // @[Mux.scala 19:72:@11053.4]
  wire [15:0] _T_5923; // @[Mux.scala 19:72:@11054.4]
  wire [15:0] _T_5938; // @[Mux.scala 19:72:@11069.4]
  wire [15:0] _T_5940; // @[Mux.scala 19:72:@11070.4]
  wire [15:0] _T_5955; // @[Mux.scala 19:72:@11085.4]
  wire [15:0] _T_5957; // @[Mux.scala 19:72:@11086.4]
  wire [15:0] _T_5958; // @[Mux.scala 19:72:@11087.4]
  wire [15:0] _T_5959; // @[Mux.scala 19:72:@11088.4]
  wire [15:0] _T_5960; // @[Mux.scala 19:72:@11089.4]
  wire [15:0] _T_5961; // @[Mux.scala 19:72:@11090.4]
  wire [15:0] _T_5962; // @[Mux.scala 19:72:@11091.4]
  wire [15:0] _T_5963; // @[Mux.scala 19:72:@11092.4]
  wire [15:0] _T_5964; // @[Mux.scala 19:72:@11093.4]
  wire [15:0] _T_5965; // @[Mux.scala 19:72:@11094.4]
  wire [15:0] _T_5966; // @[Mux.scala 19:72:@11095.4]
  wire [15:0] _T_5967; // @[Mux.scala 19:72:@11096.4]
  wire [15:0] _T_5968; // @[Mux.scala 19:72:@11097.4]
  wire [15:0] _T_5969; // @[Mux.scala 19:72:@11098.4]
  wire [15:0] _T_5970; // @[Mux.scala 19:72:@11099.4]
  wire [15:0] _T_5971; // @[Mux.scala 19:72:@11100.4]
  wire [15:0] _T_5972; // @[Mux.scala 19:72:@11101.4]
  wire  _T_6113; // @[LoadQueue.scala 121:105:@11137.4]
  wire  _T_6115; // @[LoadQueue.scala 122:18:@11138.4]
  wire  _T_6117; // @[LoadQueue.scala 122:36:@11139.4]
  wire  _T_6118; // @[LoadQueue.scala 122:27:@11140.4]
  wire  _T_6120; // @[LoadQueue.scala 122:52:@11141.4]
  wire  _T_6122; // @[LoadQueue.scala 122:85:@11142.4]
  wire  _T_6124; // @[LoadQueue.scala 122:103:@11143.4]
  wire  _T_6125; // @[LoadQueue.scala 122:94:@11144.4]
  wire  _T_6127; // @[LoadQueue.scala 122:70:@11145.4]
  wire  _T_6128; // @[LoadQueue.scala 122:67:@11146.4]
  wire  validEntriesInStoreQ_0; // @[LoadQueue.scala 121:91:@11147.4]
  wire  _T_6132; // @[LoadQueue.scala 122:18:@11149.4]
  wire  _T_6134; // @[LoadQueue.scala 122:36:@11150.4]
  wire  _T_6135; // @[LoadQueue.scala 122:27:@11151.4]
  wire  _T_6139; // @[LoadQueue.scala 122:85:@11153.4]
  wire  _T_6141; // @[LoadQueue.scala 122:103:@11154.4]
  wire  _T_6142; // @[LoadQueue.scala 122:94:@11155.4]
  wire  _T_6144; // @[LoadQueue.scala 122:70:@11156.4]
  wire  _T_6145; // @[LoadQueue.scala 122:67:@11157.4]
  wire  validEntriesInStoreQ_1; // @[LoadQueue.scala 121:91:@11158.4]
  wire  _T_6149; // @[LoadQueue.scala 122:18:@11160.4]
  wire  _T_6151; // @[LoadQueue.scala 122:36:@11161.4]
  wire  _T_6152; // @[LoadQueue.scala 122:27:@11162.4]
  wire  _T_6156; // @[LoadQueue.scala 122:85:@11164.4]
  wire  _T_6158; // @[LoadQueue.scala 122:103:@11165.4]
  wire  _T_6159; // @[LoadQueue.scala 122:94:@11166.4]
  wire  _T_6161; // @[LoadQueue.scala 122:70:@11167.4]
  wire  _T_6162; // @[LoadQueue.scala 122:67:@11168.4]
  wire  validEntriesInStoreQ_2; // @[LoadQueue.scala 121:91:@11169.4]
  wire  _T_6166; // @[LoadQueue.scala 122:18:@11171.4]
  wire  _T_6168; // @[LoadQueue.scala 122:36:@11172.4]
  wire  _T_6169; // @[LoadQueue.scala 122:27:@11173.4]
  wire  _T_6173; // @[LoadQueue.scala 122:85:@11175.4]
  wire  _T_6175; // @[LoadQueue.scala 122:103:@11176.4]
  wire  _T_6176; // @[LoadQueue.scala 122:94:@11177.4]
  wire  _T_6178; // @[LoadQueue.scala 122:70:@11178.4]
  wire  _T_6179; // @[LoadQueue.scala 122:67:@11179.4]
  wire  validEntriesInStoreQ_3; // @[LoadQueue.scala 121:91:@11180.4]
  wire  _T_6183; // @[LoadQueue.scala 122:18:@11182.4]
  wire  _T_6185; // @[LoadQueue.scala 122:36:@11183.4]
  wire  _T_6186; // @[LoadQueue.scala 122:27:@11184.4]
  wire  _T_6190; // @[LoadQueue.scala 122:85:@11186.4]
  wire  _T_6192; // @[LoadQueue.scala 122:103:@11187.4]
  wire  _T_6193; // @[LoadQueue.scala 122:94:@11188.4]
  wire  _T_6195; // @[LoadQueue.scala 122:70:@11189.4]
  wire  _T_6196; // @[LoadQueue.scala 122:67:@11190.4]
  wire  validEntriesInStoreQ_4; // @[LoadQueue.scala 121:91:@11191.4]
  wire  _T_6200; // @[LoadQueue.scala 122:18:@11193.4]
  wire  _T_6202; // @[LoadQueue.scala 122:36:@11194.4]
  wire  _T_6203; // @[LoadQueue.scala 122:27:@11195.4]
  wire  _T_6207; // @[LoadQueue.scala 122:85:@11197.4]
  wire  _T_6209; // @[LoadQueue.scala 122:103:@11198.4]
  wire  _T_6210; // @[LoadQueue.scala 122:94:@11199.4]
  wire  _T_6212; // @[LoadQueue.scala 122:70:@11200.4]
  wire  _T_6213; // @[LoadQueue.scala 122:67:@11201.4]
  wire  validEntriesInStoreQ_5; // @[LoadQueue.scala 121:91:@11202.4]
  wire  _T_6217; // @[LoadQueue.scala 122:18:@11204.4]
  wire  _T_6219; // @[LoadQueue.scala 122:36:@11205.4]
  wire  _T_6220; // @[LoadQueue.scala 122:27:@11206.4]
  wire  _T_6224; // @[LoadQueue.scala 122:85:@11208.4]
  wire  _T_6226; // @[LoadQueue.scala 122:103:@11209.4]
  wire  _T_6227; // @[LoadQueue.scala 122:94:@11210.4]
  wire  _T_6229; // @[LoadQueue.scala 122:70:@11211.4]
  wire  _T_6230; // @[LoadQueue.scala 122:67:@11212.4]
  wire  validEntriesInStoreQ_6; // @[LoadQueue.scala 121:91:@11213.4]
  wire  _T_6234; // @[LoadQueue.scala 122:18:@11215.4]
  wire  _T_6236; // @[LoadQueue.scala 122:36:@11216.4]
  wire  _T_6237; // @[LoadQueue.scala 122:27:@11217.4]
  wire  _T_6241; // @[LoadQueue.scala 122:85:@11219.4]
  wire  _T_6243; // @[LoadQueue.scala 122:103:@11220.4]
  wire  _T_6244; // @[LoadQueue.scala 122:94:@11221.4]
  wire  _T_6246; // @[LoadQueue.scala 122:70:@11222.4]
  wire  _T_6247; // @[LoadQueue.scala 122:67:@11223.4]
  wire  validEntriesInStoreQ_7; // @[LoadQueue.scala 121:91:@11224.4]
  wire  _T_6251; // @[LoadQueue.scala 122:18:@11226.4]
  wire  _T_6253; // @[LoadQueue.scala 122:36:@11227.4]
  wire  _T_6254; // @[LoadQueue.scala 122:27:@11228.4]
  wire  _T_6258; // @[LoadQueue.scala 122:85:@11230.4]
  wire  _T_6260; // @[LoadQueue.scala 122:103:@11231.4]
  wire  _T_6261; // @[LoadQueue.scala 122:94:@11232.4]
  wire  _T_6263; // @[LoadQueue.scala 122:70:@11233.4]
  wire  _T_6264; // @[LoadQueue.scala 122:67:@11234.4]
  wire  validEntriesInStoreQ_8; // @[LoadQueue.scala 121:91:@11235.4]
  wire  _T_6268; // @[LoadQueue.scala 122:18:@11237.4]
  wire  _T_6270; // @[LoadQueue.scala 122:36:@11238.4]
  wire  _T_6271; // @[LoadQueue.scala 122:27:@11239.4]
  wire  _T_6275; // @[LoadQueue.scala 122:85:@11241.4]
  wire  _T_6277; // @[LoadQueue.scala 122:103:@11242.4]
  wire  _T_6278; // @[LoadQueue.scala 122:94:@11243.4]
  wire  _T_6280; // @[LoadQueue.scala 122:70:@11244.4]
  wire  _T_6281; // @[LoadQueue.scala 122:67:@11245.4]
  wire  validEntriesInStoreQ_9; // @[LoadQueue.scala 121:91:@11246.4]
  wire  _T_6285; // @[LoadQueue.scala 122:18:@11248.4]
  wire  _T_6287; // @[LoadQueue.scala 122:36:@11249.4]
  wire  _T_6288; // @[LoadQueue.scala 122:27:@11250.4]
  wire  _T_6292; // @[LoadQueue.scala 122:85:@11252.4]
  wire  _T_6294; // @[LoadQueue.scala 122:103:@11253.4]
  wire  _T_6295; // @[LoadQueue.scala 122:94:@11254.4]
  wire  _T_6297; // @[LoadQueue.scala 122:70:@11255.4]
  wire  _T_6298; // @[LoadQueue.scala 122:67:@11256.4]
  wire  validEntriesInStoreQ_10; // @[LoadQueue.scala 121:91:@11257.4]
  wire  _T_6302; // @[LoadQueue.scala 122:18:@11259.4]
  wire  _T_6304; // @[LoadQueue.scala 122:36:@11260.4]
  wire  _T_6305; // @[LoadQueue.scala 122:27:@11261.4]
  wire  _T_6309; // @[LoadQueue.scala 122:85:@11263.4]
  wire  _T_6311; // @[LoadQueue.scala 122:103:@11264.4]
  wire  _T_6312; // @[LoadQueue.scala 122:94:@11265.4]
  wire  _T_6314; // @[LoadQueue.scala 122:70:@11266.4]
  wire  _T_6315; // @[LoadQueue.scala 122:67:@11267.4]
  wire  validEntriesInStoreQ_11; // @[LoadQueue.scala 121:91:@11268.4]
  wire  _T_6319; // @[LoadQueue.scala 122:18:@11270.4]
  wire  _T_6321; // @[LoadQueue.scala 122:36:@11271.4]
  wire  _T_6322; // @[LoadQueue.scala 122:27:@11272.4]
  wire  _T_6326; // @[LoadQueue.scala 122:85:@11274.4]
  wire  _T_6328; // @[LoadQueue.scala 122:103:@11275.4]
  wire  _T_6329; // @[LoadQueue.scala 122:94:@11276.4]
  wire  _T_6331; // @[LoadQueue.scala 122:70:@11277.4]
  wire  _T_6332; // @[LoadQueue.scala 122:67:@11278.4]
  wire  validEntriesInStoreQ_12; // @[LoadQueue.scala 121:91:@11279.4]
  wire  _T_6336; // @[LoadQueue.scala 122:18:@11281.4]
  wire  _T_6338; // @[LoadQueue.scala 122:36:@11282.4]
  wire  _T_6339; // @[LoadQueue.scala 122:27:@11283.4]
  wire  _T_6343; // @[LoadQueue.scala 122:85:@11285.4]
  wire  _T_6345; // @[LoadQueue.scala 122:103:@11286.4]
  wire  _T_6346; // @[LoadQueue.scala 122:94:@11287.4]
  wire  _T_6348; // @[LoadQueue.scala 122:70:@11288.4]
  wire  _T_6349; // @[LoadQueue.scala 122:67:@11289.4]
  wire  validEntriesInStoreQ_13; // @[LoadQueue.scala 121:91:@11290.4]
  wire  _T_6353; // @[LoadQueue.scala 122:18:@11292.4]
  wire  _T_6355; // @[LoadQueue.scala 122:36:@11293.4]
  wire  _T_6356; // @[LoadQueue.scala 122:27:@11294.4]
  wire  _T_6360; // @[LoadQueue.scala 122:85:@11296.4]
  wire  _T_6362; // @[LoadQueue.scala 122:103:@11297.4]
  wire  _T_6363; // @[LoadQueue.scala 122:94:@11298.4]
  wire  _T_6365; // @[LoadQueue.scala 122:70:@11299.4]
  wire  _T_6366; // @[LoadQueue.scala 122:67:@11300.4]
  wire  validEntriesInStoreQ_14; // @[LoadQueue.scala 121:91:@11301.4]
  wire  validEntriesInStoreQ_15; // @[LoadQueue.scala 121:91:@11312.4]
  wire  storesToCheck_0_0; // @[LoadQueue.scala 131:10:@11339.4]
  wire  _T_7654; // @[LoadQueue.scala 131:81:@11342.4]
  wire  _T_7655; // @[LoadQueue.scala 131:72:@11343.4]
  wire  _T_7657; // @[LoadQueue.scala 132:33:@11344.4]
  wire  _T_7660; // @[LoadQueue.scala 132:41:@11346.4]
  wire  _T_7662; // @[LoadQueue.scala 132:9:@11347.4]
  wire  storesToCheck_0_1; // @[LoadQueue.scala 131:10:@11348.4]
  wire  _T_7668; // @[LoadQueue.scala 131:81:@11351.4]
  wire  _T_7669; // @[LoadQueue.scala 131:72:@11352.4]
  wire  _T_7671; // @[LoadQueue.scala 132:33:@11353.4]
  wire  _T_7674; // @[LoadQueue.scala 132:41:@11355.4]
  wire  _T_7676; // @[LoadQueue.scala 132:9:@11356.4]
  wire  storesToCheck_0_2; // @[LoadQueue.scala 131:10:@11357.4]
  wire  _T_7682; // @[LoadQueue.scala 131:81:@11360.4]
  wire  _T_7683; // @[LoadQueue.scala 131:72:@11361.4]
  wire  _T_7685; // @[LoadQueue.scala 132:33:@11362.4]
  wire  _T_7688; // @[LoadQueue.scala 132:41:@11364.4]
  wire  _T_7690; // @[LoadQueue.scala 132:9:@11365.4]
  wire  storesToCheck_0_3; // @[LoadQueue.scala 131:10:@11366.4]
  wire  _T_7696; // @[LoadQueue.scala 131:81:@11369.4]
  wire  _T_7697; // @[LoadQueue.scala 131:72:@11370.4]
  wire  _T_7699; // @[LoadQueue.scala 132:33:@11371.4]
  wire  _T_7702; // @[LoadQueue.scala 132:41:@11373.4]
  wire  _T_7704; // @[LoadQueue.scala 132:9:@11374.4]
  wire  storesToCheck_0_4; // @[LoadQueue.scala 131:10:@11375.4]
  wire  _T_7710; // @[LoadQueue.scala 131:81:@11378.4]
  wire  _T_7711; // @[LoadQueue.scala 131:72:@11379.4]
  wire  _T_7713; // @[LoadQueue.scala 132:33:@11380.4]
  wire  _T_7716; // @[LoadQueue.scala 132:41:@11382.4]
  wire  _T_7718; // @[LoadQueue.scala 132:9:@11383.4]
  wire  storesToCheck_0_5; // @[LoadQueue.scala 131:10:@11384.4]
  wire  _T_7724; // @[LoadQueue.scala 131:81:@11387.4]
  wire  _T_7725; // @[LoadQueue.scala 131:72:@11388.4]
  wire  _T_7727; // @[LoadQueue.scala 132:33:@11389.4]
  wire  _T_7730; // @[LoadQueue.scala 132:41:@11391.4]
  wire  _T_7732; // @[LoadQueue.scala 132:9:@11392.4]
  wire  storesToCheck_0_6; // @[LoadQueue.scala 131:10:@11393.4]
  wire  _T_7738; // @[LoadQueue.scala 131:81:@11396.4]
  wire  _T_7739; // @[LoadQueue.scala 131:72:@11397.4]
  wire  _T_7741; // @[LoadQueue.scala 132:33:@11398.4]
  wire  _T_7744; // @[LoadQueue.scala 132:41:@11400.4]
  wire  _T_7746; // @[LoadQueue.scala 132:9:@11401.4]
  wire  storesToCheck_0_7; // @[LoadQueue.scala 131:10:@11402.4]
  wire  _T_7752; // @[LoadQueue.scala 131:81:@11405.4]
  wire  _T_7753; // @[LoadQueue.scala 131:72:@11406.4]
  wire  _T_7755; // @[LoadQueue.scala 132:33:@11407.4]
  wire  _T_7758; // @[LoadQueue.scala 132:41:@11409.4]
  wire  _T_7760; // @[LoadQueue.scala 132:9:@11410.4]
  wire  storesToCheck_0_8; // @[LoadQueue.scala 131:10:@11411.4]
  wire  _T_7766; // @[LoadQueue.scala 131:81:@11414.4]
  wire  _T_7767; // @[LoadQueue.scala 131:72:@11415.4]
  wire  _T_7769; // @[LoadQueue.scala 132:33:@11416.4]
  wire  _T_7772; // @[LoadQueue.scala 132:41:@11418.4]
  wire  _T_7774; // @[LoadQueue.scala 132:9:@11419.4]
  wire  storesToCheck_0_9; // @[LoadQueue.scala 131:10:@11420.4]
  wire  _T_7780; // @[LoadQueue.scala 131:81:@11423.4]
  wire  _T_7781; // @[LoadQueue.scala 131:72:@11424.4]
  wire  _T_7783; // @[LoadQueue.scala 132:33:@11425.4]
  wire  _T_7786; // @[LoadQueue.scala 132:41:@11427.4]
  wire  _T_7788; // @[LoadQueue.scala 132:9:@11428.4]
  wire  storesToCheck_0_10; // @[LoadQueue.scala 131:10:@11429.4]
  wire  _T_7794; // @[LoadQueue.scala 131:81:@11432.4]
  wire  _T_7795; // @[LoadQueue.scala 131:72:@11433.4]
  wire  _T_7797; // @[LoadQueue.scala 132:33:@11434.4]
  wire  _T_7800; // @[LoadQueue.scala 132:41:@11436.4]
  wire  _T_7802; // @[LoadQueue.scala 132:9:@11437.4]
  wire  storesToCheck_0_11; // @[LoadQueue.scala 131:10:@11438.4]
  wire  _T_7808; // @[LoadQueue.scala 131:81:@11441.4]
  wire  _T_7809; // @[LoadQueue.scala 131:72:@11442.4]
  wire  _T_7811; // @[LoadQueue.scala 132:33:@11443.4]
  wire  _T_7814; // @[LoadQueue.scala 132:41:@11445.4]
  wire  _T_7816; // @[LoadQueue.scala 132:9:@11446.4]
  wire  storesToCheck_0_12; // @[LoadQueue.scala 131:10:@11447.4]
  wire  _T_7822; // @[LoadQueue.scala 131:81:@11450.4]
  wire  _T_7823; // @[LoadQueue.scala 131:72:@11451.4]
  wire  _T_7825; // @[LoadQueue.scala 132:33:@11452.4]
  wire  _T_7828; // @[LoadQueue.scala 132:41:@11454.4]
  wire  _T_7830; // @[LoadQueue.scala 132:9:@11455.4]
  wire  storesToCheck_0_13; // @[LoadQueue.scala 131:10:@11456.4]
  wire  _T_7836; // @[LoadQueue.scala 131:81:@11459.4]
  wire  _T_7837; // @[LoadQueue.scala 131:72:@11460.4]
  wire  _T_7839; // @[LoadQueue.scala 132:33:@11461.4]
  wire  _T_7842; // @[LoadQueue.scala 132:41:@11463.4]
  wire  _T_7844; // @[LoadQueue.scala 132:9:@11464.4]
  wire  storesToCheck_0_14; // @[LoadQueue.scala 131:10:@11465.4]
  wire  _T_7850; // @[LoadQueue.scala 131:81:@11468.4]
  wire  storesToCheck_0_15; // @[LoadQueue.scala 131:10:@11474.4]
  wire  storesToCheck_1_0; // @[LoadQueue.scala 131:10:@11516.4]
  wire  _T_7900; // @[LoadQueue.scala 131:81:@11519.4]
  wire  _T_7901; // @[LoadQueue.scala 131:72:@11520.4]
  wire  _T_7903; // @[LoadQueue.scala 132:33:@11521.4]
  wire  _T_7906; // @[LoadQueue.scala 132:41:@11523.4]
  wire  _T_7908; // @[LoadQueue.scala 132:9:@11524.4]
  wire  storesToCheck_1_1; // @[LoadQueue.scala 131:10:@11525.4]
  wire  _T_7914; // @[LoadQueue.scala 131:81:@11528.4]
  wire  _T_7915; // @[LoadQueue.scala 131:72:@11529.4]
  wire  _T_7917; // @[LoadQueue.scala 132:33:@11530.4]
  wire  _T_7920; // @[LoadQueue.scala 132:41:@11532.4]
  wire  _T_7922; // @[LoadQueue.scala 132:9:@11533.4]
  wire  storesToCheck_1_2; // @[LoadQueue.scala 131:10:@11534.4]
  wire  _T_7928; // @[LoadQueue.scala 131:81:@11537.4]
  wire  _T_7929; // @[LoadQueue.scala 131:72:@11538.4]
  wire  _T_7931; // @[LoadQueue.scala 132:33:@11539.4]
  wire  _T_7934; // @[LoadQueue.scala 132:41:@11541.4]
  wire  _T_7936; // @[LoadQueue.scala 132:9:@11542.4]
  wire  storesToCheck_1_3; // @[LoadQueue.scala 131:10:@11543.4]
  wire  _T_7942; // @[LoadQueue.scala 131:81:@11546.4]
  wire  _T_7943; // @[LoadQueue.scala 131:72:@11547.4]
  wire  _T_7945; // @[LoadQueue.scala 132:33:@11548.4]
  wire  _T_7948; // @[LoadQueue.scala 132:41:@11550.4]
  wire  _T_7950; // @[LoadQueue.scala 132:9:@11551.4]
  wire  storesToCheck_1_4; // @[LoadQueue.scala 131:10:@11552.4]
  wire  _T_7956; // @[LoadQueue.scala 131:81:@11555.4]
  wire  _T_7957; // @[LoadQueue.scala 131:72:@11556.4]
  wire  _T_7959; // @[LoadQueue.scala 132:33:@11557.4]
  wire  _T_7962; // @[LoadQueue.scala 132:41:@11559.4]
  wire  _T_7964; // @[LoadQueue.scala 132:9:@11560.4]
  wire  storesToCheck_1_5; // @[LoadQueue.scala 131:10:@11561.4]
  wire  _T_7970; // @[LoadQueue.scala 131:81:@11564.4]
  wire  _T_7971; // @[LoadQueue.scala 131:72:@11565.4]
  wire  _T_7973; // @[LoadQueue.scala 132:33:@11566.4]
  wire  _T_7976; // @[LoadQueue.scala 132:41:@11568.4]
  wire  _T_7978; // @[LoadQueue.scala 132:9:@11569.4]
  wire  storesToCheck_1_6; // @[LoadQueue.scala 131:10:@11570.4]
  wire  _T_7984; // @[LoadQueue.scala 131:81:@11573.4]
  wire  _T_7985; // @[LoadQueue.scala 131:72:@11574.4]
  wire  _T_7987; // @[LoadQueue.scala 132:33:@11575.4]
  wire  _T_7990; // @[LoadQueue.scala 132:41:@11577.4]
  wire  _T_7992; // @[LoadQueue.scala 132:9:@11578.4]
  wire  storesToCheck_1_7; // @[LoadQueue.scala 131:10:@11579.4]
  wire  _T_7998; // @[LoadQueue.scala 131:81:@11582.4]
  wire  _T_7999; // @[LoadQueue.scala 131:72:@11583.4]
  wire  _T_8001; // @[LoadQueue.scala 132:33:@11584.4]
  wire  _T_8004; // @[LoadQueue.scala 132:41:@11586.4]
  wire  _T_8006; // @[LoadQueue.scala 132:9:@11587.4]
  wire  storesToCheck_1_8; // @[LoadQueue.scala 131:10:@11588.4]
  wire  _T_8012; // @[LoadQueue.scala 131:81:@11591.4]
  wire  _T_8013; // @[LoadQueue.scala 131:72:@11592.4]
  wire  _T_8015; // @[LoadQueue.scala 132:33:@11593.4]
  wire  _T_8018; // @[LoadQueue.scala 132:41:@11595.4]
  wire  _T_8020; // @[LoadQueue.scala 132:9:@11596.4]
  wire  storesToCheck_1_9; // @[LoadQueue.scala 131:10:@11597.4]
  wire  _T_8026; // @[LoadQueue.scala 131:81:@11600.4]
  wire  _T_8027; // @[LoadQueue.scala 131:72:@11601.4]
  wire  _T_8029; // @[LoadQueue.scala 132:33:@11602.4]
  wire  _T_8032; // @[LoadQueue.scala 132:41:@11604.4]
  wire  _T_8034; // @[LoadQueue.scala 132:9:@11605.4]
  wire  storesToCheck_1_10; // @[LoadQueue.scala 131:10:@11606.4]
  wire  _T_8040; // @[LoadQueue.scala 131:81:@11609.4]
  wire  _T_8041; // @[LoadQueue.scala 131:72:@11610.4]
  wire  _T_8043; // @[LoadQueue.scala 132:33:@11611.4]
  wire  _T_8046; // @[LoadQueue.scala 132:41:@11613.4]
  wire  _T_8048; // @[LoadQueue.scala 132:9:@11614.4]
  wire  storesToCheck_1_11; // @[LoadQueue.scala 131:10:@11615.4]
  wire  _T_8054; // @[LoadQueue.scala 131:81:@11618.4]
  wire  _T_8055; // @[LoadQueue.scala 131:72:@11619.4]
  wire  _T_8057; // @[LoadQueue.scala 132:33:@11620.4]
  wire  _T_8060; // @[LoadQueue.scala 132:41:@11622.4]
  wire  _T_8062; // @[LoadQueue.scala 132:9:@11623.4]
  wire  storesToCheck_1_12; // @[LoadQueue.scala 131:10:@11624.4]
  wire  _T_8068; // @[LoadQueue.scala 131:81:@11627.4]
  wire  _T_8069; // @[LoadQueue.scala 131:72:@11628.4]
  wire  _T_8071; // @[LoadQueue.scala 132:33:@11629.4]
  wire  _T_8074; // @[LoadQueue.scala 132:41:@11631.4]
  wire  _T_8076; // @[LoadQueue.scala 132:9:@11632.4]
  wire  storesToCheck_1_13; // @[LoadQueue.scala 131:10:@11633.4]
  wire  _T_8082; // @[LoadQueue.scala 131:81:@11636.4]
  wire  _T_8083; // @[LoadQueue.scala 131:72:@11637.4]
  wire  _T_8085; // @[LoadQueue.scala 132:33:@11638.4]
  wire  _T_8088; // @[LoadQueue.scala 132:41:@11640.4]
  wire  _T_8090; // @[LoadQueue.scala 132:9:@11641.4]
  wire  storesToCheck_1_14; // @[LoadQueue.scala 131:10:@11642.4]
  wire  _T_8096; // @[LoadQueue.scala 131:81:@11645.4]
  wire  storesToCheck_1_15; // @[LoadQueue.scala 131:10:@11651.4]
  wire  storesToCheck_2_0; // @[LoadQueue.scala 131:10:@11693.4]
  wire  _T_8146; // @[LoadQueue.scala 131:81:@11696.4]
  wire  _T_8147; // @[LoadQueue.scala 131:72:@11697.4]
  wire  _T_8149; // @[LoadQueue.scala 132:33:@11698.4]
  wire  _T_8152; // @[LoadQueue.scala 132:41:@11700.4]
  wire  _T_8154; // @[LoadQueue.scala 132:9:@11701.4]
  wire  storesToCheck_2_1; // @[LoadQueue.scala 131:10:@11702.4]
  wire  _T_8160; // @[LoadQueue.scala 131:81:@11705.4]
  wire  _T_8161; // @[LoadQueue.scala 131:72:@11706.4]
  wire  _T_8163; // @[LoadQueue.scala 132:33:@11707.4]
  wire  _T_8166; // @[LoadQueue.scala 132:41:@11709.4]
  wire  _T_8168; // @[LoadQueue.scala 132:9:@11710.4]
  wire  storesToCheck_2_2; // @[LoadQueue.scala 131:10:@11711.4]
  wire  _T_8174; // @[LoadQueue.scala 131:81:@11714.4]
  wire  _T_8175; // @[LoadQueue.scala 131:72:@11715.4]
  wire  _T_8177; // @[LoadQueue.scala 132:33:@11716.4]
  wire  _T_8180; // @[LoadQueue.scala 132:41:@11718.4]
  wire  _T_8182; // @[LoadQueue.scala 132:9:@11719.4]
  wire  storesToCheck_2_3; // @[LoadQueue.scala 131:10:@11720.4]
  wire  _T_8188; // @[LoadQueue.scala 131:81:@11723.4]
  wire  _T_8189; // @[LoadQueue.scala 131:72:@11724.4]
  wire  _T_8191; // @[LoadQueue.scala 132:33:@11725.4]
  wire  _T_8194; // @[LoadQueue.scala 132:41:@11727.4]
  wire  _T_8196; // @[LoadQueue.scala 132:9:@11728.4]
  wire  storesToCheck_2_4; // @[LoadQueue.scala 131:10:@11729.4]
  wire  _T_8202; // @[LoadQueue.scala 131:81:@11732.4]
  wire  _T_8203; // @[LoadQueue.scala 131:72:@11733.4]
  wire  _T_8205; // @[LoadQueue.scala 132:33:@11734.4]
  wire  _T_8208; // @[LoadQueue.scala 132:41:@11736.4]
  wire  _T_8210; // @[LoadQueue.scala 132:9:@11737.4]
  wire  storesToCheck_2_5; // @[LoadQueue.scala 131:10:@11738.4]
  wire  _T_8216; // @[LoadQueue.scala 131:81:@11741.4]
  wire  _T_8217; // @[LoadQueue.scala 131:72:@11742.4]
  wire  _T_8219; // @[LoadQueue.scala 132:33:@11743.4]
  wire  _T_8222; // @[LoadQueue.scala 132:41:@11745.4]
  wire  _T_8224; // @[LoadQueue.scala 132:9:@11746.4]
  wire  storesToCheck_2_6; // @[LoadQueue.scala 131:10:@11747.4]
  wire  _T_8230; // @[LoadQueue.scala 131:81:@11750.4]
  wire  _T_8231; // @[LoadQueue.scala 131:72:@11751.4]
  wire  _T_8233; // @[LoadQueue.scala 132:33:@11752.4]
  wire  _T_8236; // @[LoadQueue.scala 132:41:@11754.4]
  wire  _T_8238; // @[LoadQueue.scala 132:9:@11755.4]
  wire  storesToCheck_2_7; // @[LoadQueue.scala 131:10:@11756.4]
  wire  _T_8244; // @[LoadQueue.scala 131:81:@11759.4]
  wire  _T_8245; // @[LoadQueue.scala 131:72:@11760.4]
  wire  _T_8247; // @[LoadQueue.scala 132:33:@11761.4]
  wire  _T_8250; // @[LoadQueue.scala 132:41:@11763.4]
  wire  _T_8252; // @[LoadQueue.scala 132:9:@11764.4]
  wire  storesToCheck_2_8; // @[LoadQueue.scala 131:10:@11765.4]
  wire  _T_8258; // @[LoadQueue.scala 131:81:@11768.4]
  wire  _T_8259; // @[LoadQueue.scala 131:72:@11769.4]
  wire  _T_8261; // @[LoadQueue.scala 132:33:@11770.4]
  wire  _T_8264; // @[LoadQueue.scala 132:41:@11772.4]
  wire  _T_8266; // @[LoadQueue.scala 132:9:@11773.4]
  wire  storesToCheck_2_9; // @[LoadQueue.scala 131:10:@11774.4]
  wire  _T_8272; // @[LoadQueue.scala 131:81:@11777.4]
  wire  _T_8273; // @[LoadQueue.scala 131:72:@11778.4]
  wire  _T_8275; // @[LoadQueue.scala 132:33:@11779.4]
  wire  _T_8278; // @[LoadQueue.scala 132:41:@11781.4]
  wire  _T_8280; // @[LoadQueue.scala 132:9:@11782.4]
  wire  storesToCheck_2_10; // @[LoadQueue.scala 131:10:@11783.4]
  wire  _T_8286; // @[LoadQueue.scala 131:81:@11786.4]
  wire  _T_8287; // @[LoadQueue.scala 131:72:@11787.4]
  wire  _T_8289; // @[LoadQueue.scala 132:33:@11788.4]
  wire  _T_8292; // @[LoadQueue.scala 132:41:@11790.4]
  wire  _T_8294; // @[LoadQueue.scala 132:9:@11791.4]
  wire  storesToCheck_2_11; // @[LoadQueue.scala 131:10:@11792.4]
  wire  _T_8300; // @[LoadQueue.scala 131:81:@11795.4]
  wire  _T_8301; // @[LoadQueue.scala 131:72:@11796.4]
  wire  _T_8303; // @[LoadQueue.scala 132:33:@11797.4]
  wire  _T_8306; // @[LoadQueue.scala 132:41:@11799.4]
  wire  _T_8308; // @[LoadQueue.scala 132:9:@11800.4]
  wire  storesToCheck_2_12; // @[LoadQueue.scala 131:10:@11801.4]
  wire  _T_8314; // @[LoadQueue.scala 131:81:@11804.4]
  wire  _T_8315; // @[LoadQueue.scala 131:72:@11805.4]
  wire  _T_8317; // @[LoadQueue.scala 132:33:@11806.4]
  wire  _T_8320; // @[LoadQueue.scala 132:41:@11808.4]
  wire  _T_8322; // @[LoadQueue.scala 132:9:@11809.4]
  wire  storesToCheck_2_13; // @[LoadQueue.scala 131:10:@11810.4]
  wire  _T_8328; // @[LoadQueue.scala 131:81:@11813.4]
  wire  _T_8329; // @[LoadQueue.scala 131:72:@11814.4]
  wire  _T_8331; // @[LoadQueue.scala 132:33:@11815.4]
  wire  _T_8334; // @[LoadQueue.scala 132:41:@11817.4]
  wire  _T_8336; // @[LoadQueue.scala 132:9:@11818.4]
  wire  storesToCheck_2_14; // @[LoadQueue.scala 131:10:@11819.4]
  wire  _T_8342; // @[LoadQueue.scala 131:81:@11822.4]
  wire  storesToCheck_2_15; // @[LoadQueue.scala 131:10:@11828.4]
  wire  storesToCheck_3_0; // @[LoadQueue.scala 131:10:@11870.4]
  wire  _T_8392; // @[LoadQueue.scala 131:81:@11873.4]
  wire  _T_8393; // @[LoadQueue.scala 131:72:@11874.4]
  wire  _T_8395; // @[LoadQueue.scala 132:33:@11875.4]
  wire  _T_8398; // @[LoadQueue.scala 132:41:@11877.4]
  wire  _T_8400; // @[LoadQueue.scala 132:9:@11878.4]
  wire  storesToCheck_3_1; // @[LoadQueue.scala 131:10:@11879.4]
  wire  _T_8406; // @[LoadQueue.scala 131:81:@11882.4]
  wire  _T_8407; // @[LoadQueue.scala 131:72:@11883.4]
  wire  _T_8409; // @[LoadQueue.scala 132:33:@11884.4]
  wire  _T_8412; // @[LoadQueue.scala 132:41:@11886.4]
  wire  _T_8414; // @[LoadQueue.scala 132:9:@11887.4]
  wire  storesToCheck_3_2; // @[LoadQueue.scala 131:10:@11888.4]
  wire  _T_8420; // @[LoadQueue.scala 131:81:@11891.4]
  wire  _T_8421; // @[LoadQueue.scala 131:72:@11892.4]
  wire  _T_8423; // @[LoadQueue.scala 132:33:@11893.4]
  wire  _T_8426; // @[LoadQueue.scala 132:41:@11895.4]
  wire  _T_8428; // @[LoadQueue.scala 132:9:@11896.4]
  wire  storesToCheck_3_3; // @[LoadQueue.scala 131:10:@11897.4]
  wire  _T_8434; // @[LoadQueue.scala 131:81:@11900.4]
  wire  _T_8435; // @[LoadQueue.scala 131:72:@11901.4]
  wire  _T_8437; // @[LoadQueue.scala 132:33:@11902.4]
  wire  _T_8440; // @[LoadQueue.scala 132:41:@11904.4]
  wire  _T_8442; // @[LoadQueue.scala 132:9:@11905.4]
  wire  storesToCheck_3_4; // @[LoadQueue.scala 131:10:@11906.4]
  wire  _T_8448; // @[LoadQueue.scala 131:81:@11909.4]
  wire  _T_8449; // @[LoadQueue.scala 131:72:@11910.4]
  wire  _T_8451; // @[LoadQueue.scala 132:33:@11911.4]
  wire  _T_8454; // @[LoadQueue.scala 132:41:@11913.4]
  wire  _T_8456; // @[LoadQueue.scala 132:9:@11914.4]
  wire  storesToCheck_3_5; // @[LoadQueue.scala 131:10:@11915.4]
  wire  _T_8462; // @[LoadQueue.scala 131:81:@11918.4]
  wire  _T_8463; // @[LoadQueue.scala 131:72:@11919.4]
  wire  _T_8465; // @[LoadQueue.scala 132:33:@11920.4]
  wire  _T_8468; // @[LoadQueue.scala 132:41:@11922.4]
  wire  _T_8470; // @[LoadQueue.scala 132:9:@11923.4]
  wire  storesToCheck_3_6; // @[LoadQueue.scala 131:10:@11924.4]
  wire  _T_8476; // @[LoadQueue.scala 131:81:@11927.4]
  wire  _T_8477; // @[LoadQueue.scala 131:72:@11928.4]
  wire  _T_8479; // @[LoadQueue.scala 132:33:@11929.4]
  wire  _T_8482; // @[LoadQueue.scala 132:41:@11931.4]
  wire  _T_8484; // @[LoadQueue.scala 132:9:@11932.4]
  wire  storesToCheck_3_7; // @[LoadQueue.scala 131:10:@11933.4]
  wire  _T_8490; // @[LoadQueue.scala 131:81:@11936.4]
  wire  _T_8491; // @[LoadQueue.scala 131:72:@11937.4]
  wire  _T_8493; // @[LoadQueue.scala 132:33:@11938.4]
  wire  _T_8496; // @[LoadQueue.scala 132:41:@11940.4]
  wire  _T_8498; // @[LoadQueue.scala 132:9:@11941.4]
  wire  storesToCheck_3_8; // @[LoadQueue.scala 131:10:@11942.4]
  wire  _T_8504; // @[LoadQueue.scala 131:81:@11945.4]
  wire  _T_8505; // @[LoadQueue.scala 131:72:@11946.4]
  wire  _T_8507; // @[LoadQueue.scala 132:33:@11947.4]
  wire  _T_8510; // @[LoadQueue.scala 132:41:@11949.4]
  wire  _T_8512; // @[LoadQueue.scala 132:9:@11950.4]
  wire  storesToCheck_3_9; // @[LoadQueue.scala 131:10:@11951.4]
  wire  _T_8518; // @[LoadQueue.scala 131:81:@11954.4]
  wire  _T_8519; // @[LoadQueue.scala 131:72:@11955.4]
  wire  _T_8521; // @[LoadQueue.scala 132:33:@11956.4]
  wire  _T_8524; // @[LoadQueue.scala 132:41:@11958.4]
  wire  _T_8526; // @[LoadQueue.scala 132:9:@11959.4]
  wire  storesToCheck_3_10; // @[LoadQueue.scala 131:10:@11960.4]
  wire  _T_8532; // @[LoadQueue.scala 131:81:@11963.4]
  wire  _T_8533; // @[LoadQueue.scala 131:72:@11964.4]
  wire  _T_8535; // @[LoadQueue.scala 132:33:@11965.4]
  wire  _T_8538; // @[LoadQueue.scala 132:41:@11967.4]
  wire  _T_8540; // @[LoadQueue.scala 132:9:@11968.4]
  wire  storesToCheck_3_11; // @[LoadQueue.scala 131:10:@11969.4]
  wire  _T_8546; // @[LoadQueue.scala 131:81:@11972.4]
  wire  _T_8547; // @[LoadQueue.scala 131:72:@11973.4]
  wire  _T_8549; // @[LoadQueue.scala 132:33:@11974.4]
  wire  _T_8552; // @[LoadQueue.scala 132:41:@11976.4]
  wire  _T_8554; // @[LoadQueue.scala 132:9:@11977.4]
  wire  storesToCheck_3_12; // @[LoadQueue.scala 131:10:@11978.4]
  wire  _T_8560; // @[LoadQueue.scala 131:81:@11981.4]
  wire  _T_8561; // @[LoadQueue.scala 131:72:@11982.4]
  wire  _T_8563; // @[LoadQueue.scala 132:33:@11983.4]
  wire  _T_8566; // @[LoadQueue.scala 132:41:@11985.4]
  wire  _T_8568; // @[LoadQueue.scala 132:9:@11986.4]
  wire  storesToCheck_3_13; // @[LoadQueue.scala 131:10:@11987.4]
  wire  _T_8574; // @[LoadQueue.scala 131:81:@11990.4]
  wire  _T_8575; // @[LoadQueue.scala 131:72:@11991.4]
  wire  _T_8577; // @[LoadQueue.scala 132:33:@11992.4]
  wire  _T_8580; // @[LoadQueue.scala 132:41:@11994.4]
  wire  _T_8582; // @[LoadQueue.scala 132:9:@11995.4]
  wire  storesToCheck_3_14; // @[LoadQueue.scala 131:10:@11996.4]
  wire  _T_8588; // @[LoadQueue.scala 131:81:@11999.4]
  wire  storesToCheck_3_15; // @[LoadQueue.scala 131:10:@12005.4]
  wire  storesToCheck_4_0; // @[LoadQueue.scala 131:10:@12047.4]
  wire  _T_8638; // @[LoadQueue.scala 131:81:@12050.4]
  wire  _T_8639; // @[LoadQueue.scala 131:72:@12051.4]
  wire  _T_8641; // @[LoadQueue.scala 132:33:@12052.4]
  wire  _T_8644; // @[LoadQueue.scala 132:41:@12054.4]
  wire  _T_8646; // @[LoadQueue.scala 132:9:@12055.4]
  wire  storesToCheck_4_1; // @[LoadQueue.scala 131:10:@12056.4]
  wire  _T_8652; // @[LoadQueue.scala 131:81:@12059.4]
  wire  _T_8653; // @[LoadQueue.scala 131:72:@12060.4]
  wire  _T_8655; // @[LoadQueue.scala 132:33:@12061.4]
  wire  _T_8658; // @[LoadQueue.scala 132:41:@12063.4]
  wire  _T_8660; // @[LoadQueue.scala 132:9:@12064.4]
  wire  storesToCheck_4_2; // @[LoadQueue.scala 131:10:@12065.4]
  wire  _T_8666; // @[LoadQueue.scala 131:81:@12068.4]
  wire  _T_8667; // @[LoadQueue.scala 131:72:@12069.4]
  wire  _T_8669; // @[LoadQueue.scala 132:33:@12070.4]
  wire  _T_8672; // @[LoadQueue.scala 132:41:@12072.4]
  wire  _T_8674; // @[LoadQueue.scala 132:9:@12073.4]
  wire  storesToCheck_4_3; // @[LoadQueue.scala 131:10:@12074.4]
  wire  _T_8680; // @[LoadQueue.scala 131:81:@12077.4]
  wire  _T_8681; // @[LoadQueue.scala 131:72:@12078.4]
  wire  _T_8683; // @[LoadQueue.scala 132:33:@12079.4]
  wire  _T_8686; // @[LoadQueue.scala 132:41:@12081.4]
  wire  _T_8688; // @[LoadQueue.scala 132:9:@12082.4]
  wire  storesToCheck_4_4; // @[LoadQueue.scala 131:10:@12083.4]
  wire  _T_8694; // @[LoadQueue.scala 131:81:@12086.4]
  wire  _T_8695; // @[LoadQueue.scala 131:72:@12087.4]
  wire  _T_8697; // @[LoadQueue.scala 132:33:@12088.4]
  wire  _T_8700; // @[LoadQueue.scala 132:41:@12090.4]
  wire  _T_8702; // @[LoadQueue.scala 132:9:@12091.4]
  wire  storesToCheck_4_5; // @[LoadQueue.scala 131:10:@12092.4]
  wire  _T_8708; // @[LoadQueue.scala 131:81:@12095.4]
  wire  _T_8709; // @[LoadQueue.scala 131:72:@12096.4]
  wire  _T_8711; // @[LoadQueue.scala 132:33:@12097.4]
  wire  _T_8714; // @[LoadQueue.scala 132:41:@12099.4]
  wire  _T_8716; // @[LoadQueue.scala 132:9:@12100.4]
  wire  storesToCheck_4_6; // @[LoadQueue.scala 131:10:@12101.4]
  wire  _T_8722; // @[LoadQueue.scala 131:81:@12104.4]
  wire  _T_8723; // @[LoadQueue.scala 131:72:@12105.4]
  wire  _T_8725; // @[LoadQueue.scala 132:33:@12106.4]
  wire  _T_8728; // @[LoadQueue.scala 132:41:@12108.4]
  wire  _T_8730; // @[LoadQueue.scala 132:9:@12109.4]
  wire  storesToCheck_4_7; // @[LoadQueue.scala 131:10:@12110.4]
  wire  _T_8736; // @[LoadQueue.scala 131:81:@12113.4]
  wire  _T_8737; // @[LoadQueue.scala 131:72:@12114.4]
  wire  _T_8739; // @[LoadQueue.scala 132:33:@12115.4]
  wire  _T_8742; // @[LoadQueue.scala 132:41:@12117.4]
  wire  _T_8744; // @[LoadQueue.scala 132:9:@12118.4]
  wire  storesToCheck_4_8; // @[LoadQueue.scala 131:10:@12119.4]
  wire  _T_8750; // @[LoadQueue.scala 131:81:@12122.4]
  wire  _T_8751; // @[LoadQueue.scala 131:72:@12123.4]
  wire  _T_8753; // @[LoadQueue.scala 132:33:@12124.4]
  wire  _T_8756; // @[LoadQueue.scala 132:41:@12126.4]
  wire  _T_8758; // @[LoadQueue.scala 132:9:@12127.4]
  wire  storesToCheck_4_9; // @[LoadQueue.scala 131:10:@12128.4]
  wire  _T_8764; // @[LoadQueue.scala 131:81:@12131.4]
  wire  _T_8765; // @[LoadQueue.scala 131:72:@12132.4]
  wire  _T_8767; // @[LoadQueue.scala 132:33:@12133.4]
  wire  _T_8770; // @[LoadQueue.scala 132:41:@12135.4]
  wire  _T_8772; // @[LoadQueue.scala 132:9:@12136.4]
  wire  storesToCheck_4_10; // @[LoadQueue.scala 131:10:@12137.4]
  wire  _T_8778; // @[LoadQueue.scala 131:81:@12140.4]
  wire  _T_8779; // @[LoadQueue.scala 131:72:@12141.4]
  wire  _T_8781; // @[LoadQueue.scala 132:33:@12142.4]
  wire  _T_8784; // @[LoadQueue.scala 132:41:@12144.4]
  wire  _T_8786; // @[LoadQueue.scala 132:9:@12145.4]
  wire  storesToCheck_4_11; // @[LoadQueue.scala 131:10:@12146.4]
  wire  _T_8792; // @[LoadQueue.scala 131:81:@12149.4]
  wire  _T_8793; // @[LoadQueue.scala 131:72:@12150.4]
  wire  _T_8795; // @[LoadQueue.scala 132:33:@12151.4]
  wire  _T_8798; // @[LoadQueue.scala 132:41:@12153.4]
  wire  _T_8800; // @[LoadQueue.scala 132:9:@12154.4]
  wire  storesToCheck_4_12; // @[LoadQueue.scala 131:10:@12155.4]
  wire  _T_8806; // @[LoadQueue.scala 131:81:@12158.4]
  wire  _T_8807; // @[LoadQueue.scala 131:72:@12159.4]
  wire  _T_8809; // @[LoadQueue.scala 132:33:@12160.4]
  wire  _T_8812; // @[LoadQueue.scala 132:41:@12162.4]
  wire  _T_8814; // @[LoadQueue.scala 132:9:@12163.4]
  wire  storesToCheck_4_13; // @[LoadQueue.scala 131:10:@12164.4]
  wire  _T_8820; // @[LoadQueue.scala 131:81:@12167.4]
  wire  _T_8821; // @[LoadQueue.scala 131:72:@12168.4]
  wire  _T_8823; // @[LoadQueue.scala 132:33:@12169.4]
  wire  _T_8826; // @[LoadQueue.scala 132:41:@12171.4]
  wire  _T_8828; // @[LoadQueue.scala 132:9:@12172.4]
  wire  storesToCheck_4_14; // @[LoadQueue.scala 131:10:@12173.4]
  wire  _T_8834; // @[LoadQueue.scala 131:81:@12176.4]
  wire  storesToCheck_4_15; // @[LoadQueue.scala 131:10:@12182.4]
  wire  storesToCheck_5_0; // @[LoadQueue.scala 131:10:@12224.4]
  wire  _T_8884; // @[LoadQueue.scala 131:81:@12227.4]
  wire  _T_8885; // @[LoadQueue.scala 131:72:@12228.4]
  wire  _T_8887; // @[LoadQueue.scala 132:33:@12229.4]
  wire  _T_8890; // @[LoadQueue.scala 132:41:@12231.4]
  wire  _T_8892; // @[LoadQueue.scala 132:9:@12232.4]
  wire  storesToCheck_5_1; // @[LoadQueue.scala 131:10:@12233.4]
  wire  _T_8898; // @[LoadQueue.scala 131:81:@12236.4]
  wire  _T_8899; // @[LoadQueue.scala 131:72:@12237.4]
  wire  _T_8901; // @[LoadQueue.scala 132:33:@12238.4]
  wire  _T_8904; // @[LoadQueue.scala 132:41:@12240.4]
  wire  _T_8906; // @[LoadQueue.scala 132:9:@12241.4]
  wire  storesToCheck_5_2; // @[LoadQueue.scala 131:10:@12242.4]
  wire  _T_8912; // @[LoadQueue.scala 131:81:@12245.4]
  wire  _T_8913; // @[LoadQueue.scala 131:72:@12246.4]
  wire  _T_8915; // @[LoadQueue.scala 132:33:@12247.4]
  wire  _T_8918; // @[LoadQueue.scala 132:41:@12249.4]
  wire  _T_8920; // @[LoadQueue.scala 132:9:@12250.4]
  wire  storesToCheck_5_3; // @[LoadQueue.scala 131:10:@12251.4]
  wire  _T_8926; // @[LoadQueue.scala 131:81:@12254.4]
  wire  _T_8927; // @[LoadQueue.scala 131:72:@12255.4]
  wire  _T_8929; // @[LoadQueue.scala 132:33:@12256.4]
  wire  _T_8932; // @[LoadQueue.scala 132:41:@12258.4]
  wire  _T_8934; // @[LoadQueue.scala 132:9:@12259.4]
  wire  storesToCheck_5_4; // @[LoadQueue.scala 131:10:@12260.4]
  wire  _T_8940; // @[LoadQueue.scala 131:81:@12263.4]
  wire  _T_8941; // @[LoadQueue.scala 131:72:@12264.4]
  wire  _T_8943; // @[LoadQueue.scala 132:33:@12265.4]
  wire  _T_8946; // @[LoadQueue.scala 132:41:@12267.4]
  wire  _T_8948; // @[LoadQueue.scala 132:9:@12268.4]
  wire  storesToCheck_5_5; // @[LoadQueue.scala 131:10:@12269.4]
  wire  _T_8954; // @[LoadQueue.scala 131:81:@12272.4]
  wire  _T_8955; // @[LoadQueue.scala 131:72:@12273.4]
  wire  _T_8957; // @[LoadQueue.scala 132:33:@12274.4]
  wire  _T_8960; // @[LoadQueue.scala 132:41:@12276.4]
  wire  _T_8962; // @[LoadQueue.scala 132:9:@12277.4]
  wire  storesToCheck_5_6; // @[LoadQueue.scala 131:10:@12278.4]
  wire  _T_8968; // @[LoadQueue.scala 131:81:@12281.4]
  wire  _T_8969; // @[LoadQueue.scala 131:72:@12282.4]
  wire  _T_8971; // @[LoadQueue.scala 132:33:@12283.4]
  wire  _T_8974; // @[LoadQueue.scala 132:41:@12285.4]
  wire  _T_8976; // @[LoadQueue.scala 132:9:@12286.4]
  wire  storesToCheck_5_7; // @[LoadQueue.scala 131:10:@12287.4]
  wire  _T_8982; // @[LoadQueue.scala 131:81:@12290.4]
  wire  _T_8983; // @[LoadQueue.scala 131:72:@12291.4]
  wire  _T_8985; // @[LoadQueue.scala 132:33:@12292.4]
  wire  _T_8988; // @[LoadQueue.scala 132:41:@12294.4]
  wire  _T_8990; // @[LoadQueue.scala 132:9:@12295.4]
  wire  storesToCheck_5_8; // @[LoadQueue.scala 131:10:@12296.4]
  wire  _T_8996; // @[LoadQueue.scala 131:81:@12299.4]
  wire  _T_8997; // @[LoadQueue.scala 131:72:@12300.4]
  wire  _T_8999; // @[LoadQueue.scala 132:33:@12301.4]
  wire  _T_9002; // @[LoadQueue.scala 132:41:@12303.4]
  wire  _T_9004; // @[LoadQueue.scala 132:9:@12304.4]
  wire  storesToCheck_5_9; // @[LoadQueue.scala 131:10:@12305.4]
  wire  _T_9010; // @[LoadQueue.scala 131:81:@12308.4]
  wire  _T_9011; // @[LoadQueue.scala 131:72:@12309.4]
  wire  _T_9013; // @[LoadQueue.scala 132:33:@12310.4]
  wire  _T_9016; // @[LoadQueue.scala 132:41:@12312.4]
  wire  _T_9018; // @[LoadQueue.scala 132:9:@12313.4]
  wire  storesToCheck_5_10; // @[LoadQueue.scala 131:10:@12314.4]
  wire  _T_9024; // @[LoadQueue.scala 131:81:@12317.4]
  wire  _T_9025; // @[LoadQueue.scala 131:72:@12318.4]
  wire  _T_9027; // @[LoadQueue.scala 132:33:@12319.4]
  wire  _T_9030; // @[LoadQueue.scala 132:41:@12321.4]
  wire  _T_9032; // @[LoadQueue.scala 132:9:@12322.4]
  wire  storesToCheck_5_11; // @[LoadQueue.scala 131:10:@12323.4]
  wire  _T_9038; // @[LoadQueue.scala 131:81:@12326.4]
  wire  _T_9039; // @[LoadQueue.scala 131:72:@12327.4]
  wire  _T_9041; // @[LoadQueue.scala 132:33:@12328.4]
  wire  _T_9044; // @[LoadQueue.scala 132:41:@12330.4]
  wire  _T_9046; // @[LoadQueue.scala 132:9:@12331.4]
  wire  storesToCheck_5_12; // @[LoadQueue.scala 131:10:@12332.4]
  wire  _T_9052; // @[LoadQueue.scala 131:81:@12335.4]
  wire  _T_9053; // @[LoadQueue.scala 131:72:@12336.4]
  wire  _T_9055; // @[LoadQueue.scala 132:33:@12337.4]
  wire  _T_9058; // @[LoadQueue.scala 132:41:@12339.4]
  wire  _T_9060; // @[LoadQueue.scala 132:9:@12340.4]
  wire  storesToCheck_5_13; // @[LoadQueue.scala 131:10:@12341.4]
  wire  _T_9066; // @[LoadQueue.scala 131:81:@12344.4]
  wire  _T_9067; // @[LoadQueue.scala 131:72:@12345.4]
  wire  _T_9069; // @[LoadQueue.scala 132:33:@12346.4]
  wire  _T_9072; // @[LoadQueue.scala 132:41:@12348.4]
  wire  _T_9074; // @[LoadQueue.scala 132:9:@12349.4]
  wire  storesToCheck_5_14; // @[LoadQueue.scala 131:10:@12350.4]
  wire  _T_9080; // @[LoadQueue.scala 131:81:@12353.4]
  wire  storesToCheck_5_15; // @[LoadQueue.scala 131:10:@12359.4]
  wire  storesToCheck_6_0; // @[LoadQueue.scala 131:10:@12401.4]
  wire  _T_9130; // @[LoadQueue.scala 131:81:@12404.4]
  wire  _T_9131; // @[LoadQueue.scala 131:72:@12405.4]
  wire  _T_9133; // @[LoadQueue.scala 132:33:@12406.4]
  wire  _T_9136; // @[LoadQueue.scala 132:41:@12408.4]
  wire  _T_9138; // @[LoadQueue.scala 132:9:@12409.4]
  wire  storesToCheck_6_1; // @[LoadQueue.scala 131:10:@12410.4]
  wire  _T_9144; // @[LoadQueue.scala 131:81:@12413.4]
  wire  _T_9145; // @[LoadQueue.scala 131:72:@12414.4]
  wire  _T_9147; // @[LoadQueue.scala 132:33:@12415.4]
  wire  _T_9150; // @[LoadQueue.scala 132:41:@12417.4]
  wire  _T_9152; // @[LoadQueue.scala 132:9:@12418.4]
  wire  storesToCheck_6_2; // @[LoadQueue.scala 131:10:@12419.4]
  wire  _T_9158; // @[LoadQueue.scala 131:81:@12422.4]
  wire  _T_9159; // @[LoadQueue.scala 131:72:@12423.4]
  wire  _T_9161; // @[LoadQueue.scala 132:33:@12424.4]
  wire  _T_9164; // @[LoadQueue.scala 132:41:@12426.4]
  wire  _T_9166; // @[LoadQueue.scala 132:9:@12427.4]
  wire  storesToCheck_6_3; // @[LoadQueue.scala 131:10:@12428.4]
  wire  _T_9172; // @[LoadQueue.scala 131:81:@12431.4]
  wire  _T_9173; // @[LoadQueue.scala 131:72:@12432.4]
  wire  _T_9175; // @[LoadQueue.scala 132:33:@12433.4]
  wire  _T_9178; // @[LoadQueue.scala 132:41:@12435.4]
  wire  _T_9180; // @[LoadQueue.scala 132:9:@12436.4]
  wire  storesToCheck_6_4; // @[LoadQueue.scala 131:10:@12437.4]
  wire  _T_9186; // @[LoadQueue.scala 131:81:@12440.4]
  wire  _T_9187; // @[LoadQueue.scala 131:72:@12441.4]
  wire  _T_9189; // @[LoadQueue.scala 132:33:@12442.4]
  wire  _T_9192; // @[LoadQueue.scala 132:41:@12444.4]
  wire  _T_9194; // @[LoadQueue.scala 132:9:@12445.4]
  wire  storesToCheck_6_5; // @[LoadQueue.scala 131:10:@12446.4]
  wire  _T_9200; // @[LoadQueue.scala 131:81:@12449.4]
  wire  _T_9201; // @[LoadQueue.scala 131:72:@12450.4]
  wire  _T_9203; // @[LoadQueue.scala 132:33:@12451.4]
  wire  _T_9206; // @[LoadQueue.scala 132:41:@12453.4]
  wire  _T_9208; // @[LoadQueue.scala 132:9:@12454.4]
  wire  storesToCheck_6_6; // @[LoadQueue.scala 131:10:@12455.4]
  wire  _T_9214; // @[LoadQueue.scala 131:81:@12458.4]
  wire  _T_9215; // @[LoadQueue.scala 131:72:@12459.4]
  wire  _T_9217; // @[LoadQueue.scala 132:33:@12460.4]
  wire  _T_9220; // @[LoadQueue.scala 132:41:@12462.4]
  wire  _T_9222; // @[LoadQueue.scala 132:9:@12463.4]
  wire  storesToCheck_6_7; // @[LoadQueue.scala 131:10:@12464.4]
  wire  _T_9228; // @[LoadQueue.scala 131:81:@12467.4]
  wire  _T_9229; // @[LoadQueue.scala 131:72:@12468.4]
  wire  _T_9231; // @[LoadQueue.scala 132:33:@12469.4]
  wire  _T_9234; // @[LoadQueue.scala 132:41:@12471.4]
  wire  _T_9236; // @[LoadQueue.scala 132:9:@12472.4]
  wire  storesToCheck_6_8; // @[LoadQueue.scala 131:10:@12473.4]
  wire  _T_9242; // @[LoadQueue.scala 131:81:@12476.4]
  wire  _T_9243; // @[LoadQueue.scala 131:72:@12477.4]
  wire  _T_9245; // @[LoadQueue.scala 132:33:@12478.4]
  wire  _T_9248; // @[LoadQueue.scala 132:41:@12480.4]
  wire  _T_9250; // @[LoadQueue.scala 132:9:@12481.4]
  wire  storesToCheck_6_9; // @[LoadQueue.scala 131:10:@12482.4]
  wire  _T_9256; // @[LoadQueue.scala 131:81:@12485.4]
  wire  _T_9257; // @[LoadQueue.scala 131:72:@12486.4]
  wire  _T_9259; // @[LoadQueue.scala 132:33:@12487.4]
  wire  _T_9262; // @[LoadQueue.scala 132:41:@12489.4]
  wire  _T_9264; // @[LoadQueue.scala 132:9:@12490.4]
  wire  storesToCheck_6_10; // @[LoadQueue.scala 131:10:@12491.4]
  wire  _T_9270; // @[LoadQueue.scala 131:81:@12494.4]
  wire  _T_9271; // @[LoadQueue.scala 131:72:@12495.4]
  wire  _T_9273; // @[LoadQueue.scala 132:33:@12496.4]
  wire  _T_9276; // @[LoadQueue.scala 132:41:@12498.4]
  wire  _T_9278; // @[LoadQueue.scala 132:9:@12499.4]
  wire  storesToCheck_6_11; // @[LoadQueue.scala 131:10:@12500.4]
  wire  _T_9284; // @[LoadQueue.scala 131:81:@12503.4]
  wire  _T_9285; // @[LoadQueue.scala 131:72:@12504.4]
  wire  _T_9287; // @[LoadQueue.scala 132:33:@12505.4]
  wire  _T_9290; // @[LoadQueue.scala 132:41:@12507.4]
  wire  _T_9292; // @[LoadQueue.scala 132:9:@12508.4]
  wire  storesToCheck_6_12; // @[LoadQueue.scala 131:10:@12509.4]
  wire  _T_9298; // @[LoadQueue.scala 131:81:@12512.4]
  wire  _T_9299; // @[LoadQueue.scala 131:72:@12513.4]
  wire  _T_9301; // @[LoadQueue.scala 132:33:@12514.4]
  wire  _T_9304; // @[LoadQueue.scala 132:41:@12516.4]
  wire  _T_9306; // @[LoadQueue.scala 132:9:@12517.4]
  wire  storesToCheck_6_13; // @[LoadQueue.scala 131:10:@12518.4]
  wire  _T_9312; // @[LoadQueue.scala 131:81:@12521.4]
  wire  _T_9313; // @[LoadQueue.scala 131:72:@12522.4]
  wire  _T_9315; // @[LoadQueue.scala 132:33:@12523.4]
  wire  _T_9318; // @[LoadQueue.scala 132:41:@12525.4]
  wire  _T_9320; // @[LoadQueue.scala 132:9:@12526.4]
  wire  storesToCheck_6_14; // @[LoadQueue.scala 131:10:@12527.4]
  wire  _T_9326; // @[LoadQueue.scala 131:81:@12530.4]
  wire  storesToCheck_6_15; // @[LoadQueue.scala 131:10:@12536.4]
  wire  storesToCheck_7_0; // @[LoadQueue.scala 131:10:@12578.4]
  wire  _T_9376; // @[LoadQueue.scala 131:81:@12581.4]
  wire  _T_9377; // @[LoadQueue.scala 131:72:@12582.4]
  wire  _T_9379; // @[LoadQueue.scala 132:33:@12583.4]
  wire  _T_9382; // @[LoadQueue.scala 132:41:@12585.4]
  wire  _T_9384; // @[LoadQueue.scala 132:9:@12586.4]
  wire  storesToCheck_7_1; // @[LoadQueue.scala 131:10:@12587.4]
  wire  _T_9390; // @[LoadQueue.scala 131:81:@12590.4]
  wire  _T_9391; // @[LoadQueue.scala 131:72:@12591.4]
  wire  _T_9393; // @[LoadQueue.scala 132:33:@12592.4]
  wire  _T_9396; // @[LoadQueue.scala 132:41:@12594.4]
  wire  _T_9398; // @[LoadQueue.scala 132:9:@12595.4]
  wire  storesToCheck_7_2; // @[LoadQueue.scala 131:10:@12596.4]
  wire  _T_9404; // @[LoadQueue.scala 131:81:@12599.4]
  wire  _T_9405; // @[LoadQueue.scala 131:72:@12600.4]
  wire  _T_9407; // @[LoadQueue.scala 132:33:@12601.4]
  wire  _T_9410; // @[LoadQueue.scala 132:41:@12603.4]
  wire  _T_9412; // @[LoadQueue.scala 132:9:@12604.4]
  wire  storesToCheck_7_3; // @[LoadQueue.scala 131:10:@12605.4]
  wire  _T_9418; // @[LoadQueue.scala 131:81:@12608.4]
  wire  _T_9419; // @[LoadQueue.scala 131:72:@12609.4]
  wire  _T_9421; // @[LoadQueue.scala 132:33:@12610.4]
  wire  _T_9424; // @[LoadQueue.scala 132:41:@12612.4]
  wire  _T_9426; // @[LoadQueue.scala 132:9:@12613.4]
  wire  storesToCheck_7_4; // @[LoadQueue.scala 131:10:@12614.4]
  wire  _T_9432; // @[LoadQueue.scala 131:81:@12617.4]
  wire  _T_9433; // @[LoadQueue.scala 131:72:@12618.4]
  wire  _T_9435; // @[LoadQueue.scala 132:33:@12619.4]
  wire  _T_9438; // @[LoadQueue.scala 132:41:@12621.4]
  wire  _T_9440; // @[LoadQueue.scala 132:9:@12622.4]
  wire  storesToCheck_7_5; // @[LoadQueue.scala 131:10:@12623.4]
  wire  _T_9446; // @[LoadQueue.scala 131:81:@12626.4]
  wire  _T_9447; // @[LoadQueue.scala 131:72:@12627.4]
  wire  _T_9449; // @[LoadQueue.scala 132:33:@12628.4]
  wire  _T_9452; // @[LoadQueue.scala 132:41:@12630.4]
  wire  _T_9454; // @[LoadQueue.scala 132:9:@12631.4]
  wire  storesToCheck_7_6; // @[LoadQueue.scala 131:10:@12632.4]
  wire  _T_9460; // @[LoadQueue.scala 131:81:@12635.4]
  wire  _T_9461; // @[LoadQueue.scala 131:72:@12636.4]
  wire  _T_9463; // @[LoadQueue.scala 132:33:@12637.4]
  wire  _T_9466; // @[LoadQueue.scala 132:41:@12639.4]
  wire  _T_9468; // @[LoadQueue.scala 132:9:@12640.4]
  wire  storesToCheck_7_7; // @[LoadQueue.scala 131:10:@12641.4]
  wire  _T_9474; // @[LoadQueue.scala 131:81:@12644.4]
  wire  _T_9475; // @[LoadQueue.scala 131:72:@12645.4]
  wire  _T_9477; // @[LoadQueue.scala 132:33:@12646.4]
  wire  _T_9480; // @[LoadQueue.scala 132:41:@12648.4]
  wire  _T_9482; // @[LoadQueue.scala 132:9:@12649.4]
  wire  storesToCheck_7_8; // @[LoadQueue.scala 131:10:@12650.4]
  wire  _T_9488; // @[LoadQueue.scala 131:81:@12653.4]
  wire  _T_9489; // @[LoadQueue.scala 131:72:@12654.4]
  wire  _T_9491; // @[LoadQueue.scala 132:33:@12655.4]
  wire  _T_9494; // @[LoadQueue.scala 132:41:@12657.4]
  wire  _T_9496; // @[LoadQueue.scala 132:9:@12658.4]
  wire  storesToCheck_7_9; // @[LoadQueue.scala 131:10:@12659.4]
  wire  _T_9502; // @[LoadQueue.scala 131:81:@12662.4]
  wire  _T_9503; // @[LoadQueue.scala 131:72:@12663.4]
  wire  _T_9505; // @[LoadQueue.scala 132:33:@12664.4]
  wire  _T_9508; // @[LoadQueue.scala 132:41:@12666.4]
  wire  _T_9510; // @[LoadQueue.scala 132:9:@12667.4]
  wire  storesToCheck_7_10; // @[LoadQueue.scala 131:10:@12668.4]
  wire  _T_9516; // @[LoadQueue.scala 131:81:@12671.4]
  wire  _T_9517; // @[LoadQueue.scala 131:72:@12672.4]
  wire  _T_9519; // @[LoadQueue.scala 132:33:@12673.4]
  wire  _T_9522; // @[LoadQueue.scala 132:41:@12675.4]
  wire  _T_9524; // @[LoadQueue.scala 132:9:@12676.4]
  wire  storesToCheck_7_11; // @[LoadQueue.scala 131:10:@12677.4]
  wire  _T_9530; // @[LoadQueue.scala 131:81:@12680.4]
  wire  _T_9531; // @[LoadQueue.scala 131:72:@12681.4]
  wire  _T_9533; // @[LoadQueue.scala 132:33:@12682.4]
  wire  _T_9536; // @[LoadQueue.scala 132:41:@12684.4]
  wire  _T_9538; // @[LoadQueue.scala 132:9:@12685.4]
  wire  storesToCheck_7_12; // @[LoadQueue.scala 131:10:@12686.4]
  wire  _T_9544; // @[LoadQueue.scala 131:81:@12689.4]
  wire  _T_9545; // @[LoadQueue.scala 131:72:@12690.4]
  wire  _T_9547; // @[LoadQueue.scala 132:33:@12691.4]
  wire  _T_9550; // @[LoadQueue.scala 132:41:@12693.4]
  wire  _T_9552; // @[LoadQueue.scala 132:9:@12694.4]
  wire  storesToCheck_7_13; // @[LoadQueue.scala 131:10:@12695.4]
  wire  _T_9558; // @[LoadQueue.scala 131:81:@12698.4]
  wire  _T_9559; // @[LoadQueue.scala 131:72:@12699.4]
  wire  _T_9561; // @[LoadQueue.scala 132:33:@12700.4]
  wire  _T_9564; // @[LoadQueue.scala 132:41:@12702.4]
  wire  _T_9566; // @[LoadQueue.scala 132:9:@12703.4]
  wire  storesToCheck_7_14; // @[LoadQueue.scala 131:10:@12704.4]
  wire  _T_9572; // @[LoadQueue.scala 131:81:@12707.4]
  wire  storesToCheck_7_15; // @[LoadQueue.scala 131:10:@12713.4]
  wire  storesToCheck_8_0; // @[LoadQueue.scala 131:10:@12755.4]
  wire  _T_9622; // @[LoadQueue.scala 131:81:@12758.4]
  wire  _T_9623; // @[LoadQueue.scala 131:72:@12759.4]
  wire  _T_9625; // @[LoadQueue.scala 132:33:@12760.4]
  wire  _T_9628; // @[LoadQueue.scala 132:41:@12762.4]
  wire  _T_9630; // @[LoadQueue.scala 132:9:@12763.4]
  wire  storesToCheck_8_1; // @[LoadQueue.scala 131:10:@12764.4]
  wire  _T_9636; // @[LoadQueue.scala 131:81:@12767.4]
  wire  _T_9637; // @[LoadQueue.scala 131:72:@12768.4]
  wire  _T_9639; // @[LoadQueue.scala 132:33:@12769.4]
  wire  _T_9642; // @[LoadQueue.scala 132:41:@12771.4]
  wire  _T_9644; // @[LoadQueue.scala 132:9:@12772.4]
  wire  storesToCheck_8_2; // @[LoadQueue.scala 131:10:@12773.4]
  wire  _T_9650; // @[LoadQueue.scala 131:81:@12776.4]
  wire  _T_9651; // @[LoadQueue.scala 131:72:@12777.4]
  wire  _T_9653; // @[LoadQueue.scala 132:33:@12778.4]
  wire  _T_9656; // @[LoadQueue.scala 132:41:@12780.4]
  wire  _T_9658; // @[LoadQueue.scala 132:9:@12781.4]
  wire  storesToCheck_8_3; // @[LoadQueue.scala 131:10:@12782.4]
  wire  _T_9664; // @[LoadQueue.scala 131:81:@12785.4]
  wire  _T_9665; // @[LoadQueue.scala 131:72:@12786.4]
  wire  _T_9667; // @[LoadQueue.scala 132:33:@12787.4]
  wire  _T_9670; // @[LoadQueue.scala 132:41:@12789.4]
  wire  _T_9672; // @[LoadQueue.scala 132:9:@12790.4]
  wire  storesToCheck_8_4; // @[LoadQueue.scala 131:10:@12791.4]
  wire  _T_9678; // @[LoadQueue.scala 131:81:@12794.4]
  wire  _T_9679; // @[LoadQueue.scala 131:72:@12795.4]
  wire  _T_9681; // @[LoadQueue.scala 132:33:@12796.4]
  wire  _T_9684; // @[LoadQueue.scala 132:41:@12798.4]
  wire  _T_9686; // @[LoadQueue.scala 132:9:@12799.4]
  wire  storesToCheck_8_5; // @[LoadQueue.scala 131:10:@12800.4]
  wire  _T_9692; // @[LoadQueue.scala 131:81:@12803.4]
  wire  _T_9693; // @[LoadQueue.scala 131:72:@12804.4]
  wire  _T_9695; // @[LoadQueue.scala 132:33:@12805.4]
  wire  _T_9698; // @[LoadQueue.scala 132:41:@12807.4]
  wire  _T_9700; // @[LoadQueue.scala 132:9:@12808.4]
  wire  storesToCheck_8_6; // @[LoadQueue.scala 131:10:@12809.4]
  wire  _T_9706; // @[LoadQueue.scala 131:81:@12812.4]
  wire  _T_9707; // @[LoadQueue.scala 131:72:@12813.4]
  wire  _T_9709; // @[LoadQueue.scala 132:33:@12814.4]
  wire  _T_9712; // @[LoadQueue.scala 132:41:@12816.4]
  wire  _T_9714; // @[LoadQueue.scala 132:9:@12817.4]
  wire  storesToCheck_8_7; // @[LoadQueue.scala 131:10:@12818.4]
  wire  _T_9720; // @[LoadQueue.scala 131:81:@12821.4]
  wire  _T_9721; // @[LoadQueue.scala 131:72:@12822.4]
  wire  _T_9723; // @[LoadQueue.scala 132:33:@12823.4]
  wire  _T_9726; // @[LoadQueue.scala 132:41:@12825.4]
  wire  _T_9728; // @[LoadQueue.scala 132:9:@12826.4]
  wire  storesToCheck_8_8; // @[LoadQueue.scala 131:10:@12827.4]
  wire  _T_9734; // @[LoadQueue.scala 131:81:@12830.4]
  wire  _T_9735; // @[LoadQueue.scala 131:72:@12831.4]
  wire  _T_9737; // @[LoadQueue.scala 132:33:@12832.4]
  wire  _T_9740; // @[LoadQueue.scala 132:41:@12834.4]
  wire  _T_9742; // @[LoadQueue.scala 132:9:@12835.4]
  wire  storesToCheck_8_9; // @[LoadQueue.scala 131:10:@12836.4]
  wire  _T_9748; // @[LoadQueue.scala 131:81:@12839.4]
  wire  _T_9749; // @[LoadQueue.scala 131:72:@12840.4]
  wire  _T_9751; // @[LoadQueue.scala 132:33:@12841.4]
  wire  _T_9754; // @[LoadQueue.scala 132:41:@12843.4]
  wire  _T_9756; // @[LoadQueue.scala 132:9:@12844.4]
  wire  storesToCheck_8_10; // @[LoadQueue.scala 131:10:@12845.4]
  wire  _T_9762; // @[LoadQueue.scala 131:81:@12848.4]
  wire  _T_9763; // @[LoadQueue.scala 131:72:@12849.4]
  wire  _T_9765; // @[LoadQueue.scala 132:33:@12850.4]
  wire  _T_9768; // @[LoadQueue.scala 132:41:@12852.4]
  wire  _T_9770; // @[LoadQueue.scala 132:9:@12853.4]
  wire  storesToCheck_8_11; // @[LoadQueue.scala 131:10:@12854.4]
  wire  _T_9776; // @[LoadQueue.scala 131:81:@12857.4]
  wire  _T_9777; // @[LoadQueue.scala 131:72:@12858.4]
  wire  _T_9779; // @[LoadQueue.scala 132:33:@12859.4]
  wire  _T_9782; // @[LoadQueue.scala 132:41:@12861.4]
  wire  _T_9784; // @[LoadQueue.scala 132:9:@12862.4]
  wire  storesToCheck_8_12; // @[LoadQueue.scala 131:10:@12863.4]
  wire  _T_9790; // @[LoadQueue.scala 131:81:@12866.4]
  wire  _T_9791; // @[LoadQueue.scala 131:72:@12867.4]
  wire  _T_9793; // @[LoadQueue.scala 132:33:@12868.4]
  wire  _T_9796; // @[LoadQueue.scala 132:41:@12870.4]
  wire  _T_9798; // @[LoadQueue.scala 132:9:@12871.4]
  wire  storesToCheck_8_13; // @[LoadQueue.scala 131:10:@12872.4]
  wire  _T_9804; // @[LoadQueue.scala 131:81:@12875.4]
  wire  _T_9805; // @[LoadQueue.scala 131:72:@12876.4]
  wire  _T_9807; // @[LoadQueue.scala 132:33:@12877.4]
  wire  _T_9810; // @[LoadQueue.scala 132:41:@12879.4]
  wire  _T_9812; // @[LoadQueue.scala 132:9:@12880.4]
  wire  storesToCheck_8_14; // @[LoadQueue.scala 131:10:@12881.4]
  wire  _T_9818; // @[LoadQueue.scala 131:81:@12884.4]
  wire  storesToCheck_8_15; // @[LoadQueue.scala 131:10:@12890.4]
  wire  storesToCheck_9_0; // @[LoadQueue.scala 131:10:@12932.4]
  wire  _T_9868; // @[LoadQueue.scala 131:81:@12935.4]
  wire  _T_9869; // @[LoadQueue.scala 131:72:@12936.4]
  wire  _T_9871; // @[LoadQueue.scala 132:33:@12937.4]
  wire  _T_9874; // @[LoadQueue.scala 132:41:@12939.4]
  wire  _T_9876; // @[LoadQueue.scala 132:9:@12940.4]
  wire  storesToCheck_9_1; // @[LoadQueue.scala 131:10:@12941.4]
  wire  _T_9882; // @[LoadQueue.scala 131:81:@12944.4]
  wire  _T_9883; // @[LoadQueue.scala 131:72:@12945.4]
  wire  _T_9885; // @[LoadQueue.scala 132:33:@12946.4]
  wire  _T_9888; // @[LoadQueue.scala 132:41:@12948.4]
  wire  _T_9890; // @[LoadQueue.scala 132:9:@12949.4]
  wire  storesToCheck_9_2; // @[LoadQueue.scala 131:10:@12950.4]
  wire  _T_9896; // @[LoadQueue.scala 131:81:@12953.4]
  wire  _T_9897; // @[LoadQueue.scala 131:72:@12954.4]
  wire  _T_9899; // @[LoadQueue.scala 132:33:@12955.4]
  wire  _T_9902; // @[LoadQueue.scala 132:41:@12957.4]
  wire  _T_9904; // @[LoadQueue.scala 132:9:@12958.4]
  wire  storesToCheck_9_3; // @[LoadQueue.scala 131:10:@12959.4]
  wire  _T_9910; // @[LoadQueue.scala 131:81:@12962.4]
  wire  _T_9911; // @[LoadQueue.scala 131:72:@12963.4]
  wire  _T_9913; // @[LoadQueue.scala 132:33:@12964.4]
  wire  _T_9916; // @[LoadQueue.scala 132:41:@12966.4]
  wire  _T_9918; // @[LoadQueue.scala 132:9:@12967.4]
  wire  storesToCheck_9_4; // @[LoadQueue.scala 131:10:@12968.4]
  wire  _T_9924; // @[LoadQueue.scala 131:81:@12971.4]
  wire  _T_9925; // @[LoadQueue.scala 131:72:@12972.4]
  wire  _T_9927; // @[LoadQueue.scala 132:33:@12973.4]
  wire  _T_9930; // @[LoadQueue.scala 132:41:@12975.4]
  wire  _T_9932; // @[LoadQueue.scala 132:9:@12976.4]
  wire  storesToCheck_9_5; // @[LoadQueue.scala 131:10:@12977.4]
  wire  _T_9938; // @[LoadQueue.scala 131:81:@12980.4]
  wire  _T_9939; // @[LoadQueue.scala 131:72:@12981.4]
  wire  _T_9941; // @[LoadQueue.scala 132:33:@12982.4]
  wire  _T_9944; // @[LoadQueue.scala 132:41:@12984.4]
  wire  _T_9946; // @[LoadQueue.scala 132:9:@12985.4]
  wire  storesToCheck_9_6; // @[LoadQueue.scala 131:10:@12986.4]
  wire  _T_9952; // @[LoadQueue.scala 131:81:@12989.4]
  wire  _T_9953; // @[LoadQueue.scala 131:72:@12990.4]
  wire  _T_9955; // @[LoadQueue.scala 132:33:@12991.4]
  wire  _T_9958; // @[LoadQueue.scala 132:41:@12993.4]
  wire  _T_9960; // @[LoadQueue.scala 132:9:@12994.4]
  wire  storesToCheck_9_7; // @[LoadQueue.scala 131:10:@12995.4]
  wire  _T_9966; // @[LoadQueue.scala 131:81:@12998.4]
  wire  _T_9967; // @[LoadQueue.scala 131:72:@12999.4]
  wire  _T_9969; // @[LoadQueue.scala 132:33:@13000.4]
  wire  _T_9972; // @[LoadQueue.scala 132:41:@13002.4]
  wire  _T_9974; // @[LoadQueue.scala 132:9:@13003.4]
  wire  storesToCheck_9_8; // @[LoadQueue.scala 131:10:@13004.4]
  wire  _T_9980; // @[LoadQueue.scala 131:81:@13007.4]
  wire  _T_9981; // @[LoadQueue.scala 131:72:@13008.4]
  wire  _T_9983; // @[LoadQueue.scala 132:33:@13009.4]
  wire  _T_9986; // @[LoadQueue.scala 132:41:@13011.4]
  wire  _T_9988; // @[LoadQueue.scala 132:9:@13012.4]
  wire  storesToCheck_9_9; // @[LoadQueue.scala 131:10:@13013.4]
  wire  _T_9994; // @[LoadQueue.scala 131:81:@13016.4]
  wire  _T_9995; // @[LoadQueue.scala 131:72:@13017.4]
  wire  _T_9997; // @[LoadQueue.scala 132:33:@13018.4]
  wire  _T_10000; // @[LoadQueue.scala 132:41:@13020.4]
  wire  _T_10002; // @[LoadQueue.scala 132:9:@13021.4]
  wire  storesToCheck_9_10; // @[LoadQueue.scala 131:10:@13022.4]
  wire  _T_10008; // @[LoadQueue.scala 131:81:@13025.4]
  wire  _T_10009; // @[LoadQueue.scala 131:72:@13026.4]
  wire  _T_10011; // @[LoadQueue.scala 132:33:@13027.4]
  wire  _T_10014; // @[LoadQueue.scala 132:41:@13029.4]
  wire  _T_10016; // @[LoadQueue.scala 132:9:@13030.4]
  wire  storesToCheck_9_11; // @[LoadQueue.scala 131:10:@13031.4]
  wire  _T_10022; // @[LoadQueue.scala 131:81:@13034.4]
  wire  _T_10023; // @[LoadQueue.scala 131:72:@13035.4]
  wire  _T_10025; // @[LoadQueue.scala 132:33:@13036.4]
  wire  _T_10028; // @[LoadQueue.scala 132:41:@13038.4]
  wire  _T_10030; // @[LoadQueue.scala 132:9:@13039.4]
  wire  storesToCheck_9_12; // @[LoadQueue.scala 131:10:@13040.4]
  wire  _T_10036; // @[LoadQueue.scala 131:81:@13043.4]
  wire  _T_10037; // @[LoadQueue.scala 131:72:@13044.4]
  wire  _T_10039; // @[LoadQueue.scala 132:33:@13045.4]
  wire  _T_10042; // @[LoadQueue.scala 132:41:@13047.4]
  wire  _T_10044; // @[LoadQueue.scala 132:9:@13048.4]
  wire  storesToCheck_9_13; // @[LoadQueue.scala 131:10:@13049.4]
  wire  _T_10050; // @[LoadQueue.scala 131:81:@13052.4]
  wire  _T_10051; // @[LoadQueue.scala 131:72:@13053.4]
  wire  _T_10053; // @[LoadQueue.scala 132:33:@13054.4]
  wire  _T_10056; // @[LoadQueue.scala 132:41:@13056.4]
  wire  _T_10058; // @[LoadQueue.scala 132:9:@13057.4]
  wire  storesToCheck_9_14; // @[LoadQueue.scala 131:10:@13058.4]
  wire  _T_10064; // @[LoadQueue.scala 131:81:@13061.4]
  wire  storesToCheck_9_15; // @[LoadQueue.scala 131:10:@13067.4]
  wire  storesToCheck_10_0; // @[LoadQueue.scala 131:10:@13109.4]
  wire  _T_10114; // @[LoadQueue.scala 131:81:@13112.4]
  wire  _T_10115; // @[LoadQueue.scala 131:72:@13113.4]
  wire  _T_10117; // @[LoadQueue.scala 132:33:@13114.4]
  wire  _T_10120; // @[LoadQueue.scala 132:41:@13116.4]
  wire  _T_10122; // @[LoadQueue.scala 132:9:@13117.4]
  wire  storesToCheck_10_1; // @[LoadQueue.scala 131:10:@13118.4]
  wire  _T_10128; // @[LoadQueue.scala 131:81:@13121.4]
  wire  _T_10129; // @[LoadQueue.scala 131:72:@13122.4]
  wire  _T_10131; // @[LoadQueue.scala 132:33:@13123.4]
  wire  _T_10134; // @[LoadQueue.scala 132:41:@13125.4]
  wire  _T_10136; // @[LoadQueue.scala 132:9:@13126.4]
  wire  storesToCheck_10_2; // @[LoadQueue.scala 131:10:@13127.4]
  wire  _T_10142; // @[LoadQueue.scala 131:81:@13130.4]
  wire  _T_10143; // @[LoadQueue.scala 131:72:@13131.4]
  wire  _T_10145; // @[LoadQueue.scala 132:33:@13132.4]
  wire  _T_10148; // @[LoadQueue.scala 132:41:@13134.4]
  wire  _T_10150; // @[LoadQueue.scala 132:9:@13135.4]
  wire  storesToCheck_10_3; // @[LoadQueue.scala 131:10:@13136.4]
  wire  _T_10156; // @[LoadQueue.scala 131:81:@13139.4]
  wire  _T_10157; // @[LoadQueue.scala 131:72:@13140.4]
  wire  _T_10159; // @[LoadQueue.scala 132:33:@13141.4]
  wire  _T_10162; // @[LoadQueue.scala 132:41:@13143.4]
  wire  _T_10164; // @[LoadQueue.scala 132:9:@13144.4]
  wire  storesToCheck_10_4; // @[LoadQueue.scala 131:10:@13145.4]
  wire  _T_10170; // @[LoadQueue.scala 131:81:@13148.4]
  wire  _T_10171; // @[LoadQueue.scala 131:72:@13149.4]
  wire  _T_10173; // @[LoadQueue.scala 132:33:@13150.4]
  wire  _T_10176; // @[LoadQueue.scala 132:41:@13152.4]
  wire  _T_10178; // @[LoadQueue.scala 132:9:@13153.4]
  wire  storesToCheck_10_5; // @[LoadQueue.scala 131:10:@13154.4]
  wire  _T_10184; // @[LoadQueue.scala 131:81:@13157.4]
  wire  _T_10185; // @[LoadQueue.scala 131:72:@13158.4]
  wire  _T_10187; // @[LoadQueue.scala 132:33:@13159.4]
  wire  _T_10190; // @[LoadQueue.scala 132:41:@13161.4]
  wire  _T_10192; // @[LoadQueue.scala 132:9:@13162.4]
  wire  storesToCheck_10_6; // @[LoadQueue.scala 131:10:@13163.4]
  wire  _T_10198; // @[LoadQueue.scala 131:81:@13166.4]
  wire  _T_10199; // @[LoadQueue.scala 131:72:@13167.4]
  wire  _T_10201; // @[LoadQueue.scala 132:33:@13168.4]
  wire  _T_10204; // @[LoadQueue.scala 132:41:@13170.4]
  wire  _T_10206; // @[LoadQueue.scala 132:9:@13171.4]
  wire  storesToCheck_10_7; // @[LoadQueue.scala 131:10:@13172.4]
  wire  _T_10212; // @[LoadQueue.scala 131:81:@13175.4]
  wire  _T_10213; // @[LoadQueue.scala 131:72:@13176.4]
  wire  _T_10215; // @[LoadQueue.scala 132:33:@13177.4]
  wire  _T_10218; // @[LoadQueue.scala 132:41:@13179.4]
  wire  _T_10220; // @[LoadQueue.scala 132:9:@13180.4]
  wire  storesToCheck_10_8; // @[LoadQueue.scala 131:10:@13181.4]
  wire  _T_10226; // @[LoadQueue.scala 131:81:@13184.4]
  wire  _T_10227; // @[LoadQueue.scala 131:72:@13185.4]
  wire  _T_10229; // @[LoadQueue.scala 132:33:@13186.4]
  wire  _T_10232; // @[LoadQueue.scala 132:41:@13188.4]
  wire  _T_10234; // @[LoadQueue.scala 132:9:@13189.4]
  wire  storesToCheck_10_9; // @[LoadQueue.scala 131:10:@13190.4]
  wire  _T_10240; // @[LoadQueue.scala 131:81:@13193.4]
  wire  _T_10241; // @[LoadQueue.scala 131:72:@13194.4]
  wire  _T_10243; // @[LoadQueue.scala 132:33:@13195.4]
  wire  _T_10246; // @[LoadQueue.scala 132:41:@13197.4]
  wire  _T_10248; // @[LoadQueue.scala 132:9:@13198.4]
  wire  storesToCheck_10_10; // @[LoadQueue.scala 131:10:@13199.4]
  wire  _T_10254; // @[LoadQueue.scala 131:81:@13202.4]
  wire  _T_10255; // @[LoadQueue.scala 131:72:@13203.4]
  wire  _T_10257; // @[LoadQueue.scala 132:33:@13204.4]
  wire  _T_10260; // @[LoadQueue.scala 132:41:@13206.4]
  wire  _T_10262; // @[LoadQueue.scala 132:9:@13207.4]
  wire  storesToCheck_10_11; // @[LoadQueue.scala 131:10:@13208.4]
  wire  _T_10268; // @[LoadQueue.scala 131:81:@13211.4]
  wire  _T_10269; // @[LoadQueue.scala 131:72:@13212.4]
  wire  _T_10271; // @[LoadQueue.scala 132:33:@13213.4]
  wire  _T_10274; // @[LoadQueue.scala 132:41:@13215.4]
  wire  _T_10276; // @[LoadQueue.scala 132:9:@13216.4]
  wire  storesToCheck_10_12; // @[LoadQueue.scala 131:10:@13217.4]
  wire  _T_10282; // @[LoadQueue.scala 131:81:@13220.4]
  wire  _T_10283; // @[LoadQueue.scala 131:72:@13221.4]
  wire  _T_10285; // @[LoadQueue.scala 132:33:@13222.4]
  wire  _T_10288; // @[LoadQueue.scala 132:41:@13224.4]
  wire  _T_10290; // @[LoadQueue.scala 132:9:@13225.4]
  wire  storesToCheck_10_13; // @[LoadQueue.scala 131:10:@13226.4]
  wire  _T_10296; // @[LoadQueue.scala 131:81:@13229.4]
  wire  _T_10297; // @[LoadQueue.scala 131:72:@13230.4]
  wire  _T_10299; // @[LoadQueue.scala 132:33:@13231.4]
  wire  _T_10302; // @[LoadQueue.scala 132:41:@13233.4]
  wire  _T_10304; // @[LoadQueue.scala 132:9:@13234.4]
  wire  storesToCheck_10_14; // @[LoadQueue.scala 131:10:@13235.4]
  wire  _T_10310; // @[LoadQueue.scala 131:81:@13238.4]
  wire  storesToCheck_10_15; // @[LoadQueue.scala 131:10:@13244.4]
  wire  storesToCheck_11_0; // @[LoadQueue.scala 131:10:@13286.4]
  wire  _T_10360; // @[LoadQueue.scala 131:81:@13289.4]
  wire  _T_10361; // @[LoadQueue.scala 131:72:@13290.4]
  wire  _T_10363; // @[LoadQueue.scala 132:33:@13291.4]
  wire  _T_10366; // @[LoadQueue.scala 132:41:@13293.4]
  wire  _T_10368; // @[LoadQueue.scala 132:9:@13294.4]
  wire  storesToCheck_11_1; // @[LoadQueue.scala 131:10:@13295.4]
  wire  _T_10374; // @[LoadQueue.scala 131:81:@13298.4]
  wire  _T_10375; // @[LoadQueue.scala 131:72:@13299.4]
  wire  _T_10377; // @[LoadQueue.scala 132:33:@13300.4]
  wire  _T_10380; // @[LoadQueue.scala 132:41:@13302.4]
  wire  _T_10382; // @[LoadQueue.scala 132:9:@13303.4]
  wire  storesToCheck_11_2; // @[LoadQueue.scala 131:10:@13304.4]
  wire  _T_10388; // @[LoadQueue.scala 131:81:@13307.4]
  wire  _T_10389; // @[LoadQueue.scala 131:72:@13308.4]
  wire  _T_10391; // @[LoadQueue.scala 132:33:@13309.4]
  wire  _T_10394; // @[LoadQueue.scala 132:41:@13311.4]
  wire  _T_10396; // @[LoadQueue.scala 132:9:@13312.4]
  wire  storesToCheck_11_3; // @[LoadQueue.scala 131:10:@13313.4]
  wire  _T_10402; // @[LoadQueue.scala 131:81:@13316.4]
  wire  _T_10403; // @[LoadQueue.scala 131:72:@13317.4]
  wire  _T_10405; // @[LoadQueue.scala 132:33:@13318.4]
  wire  _T_10408; // @[LoadQueue.scala 132:41:@13320.4]
  wire  _T_10410; // @[LoadQueue.scala 132:9:@13321.4]
  wire  storesToCheck_11_4; // @[LoadQueue.scala 131:10:@13322.4]
  wire  _T_10416; // @[LoadQueue.scala 131:81:@13325.4]
  wire  _T_10417; // @[LoadQueue.scala 131:72:@13326.4]
  wire  _T_10419; // @[LoadQueue.scala 132:33:@13327.4]
  wire  _T_10422; // @[LoadQueue.scala 132:41:@13329.4]
  wire  _T_10424; // @[LoadQueue.scala 132:9:@13330.4]
  wire  storesToCheck_11_5; // @[LoadQueue.scala 131:10:@13331.4]
  wire  _T_10430; // @[LoadQueue.scala 131:81:@13334.4]
  wire  _T_10431; // @[LoadQueue.scala 131:72:@13335.4]
  wire  _T_10433; // @[LoadQueue.scala 132:33:@13336.4]
  wire  _T_10436; // @[LoadQueue.scala 132:41:@13338.4]
  wire  _T_10438; // @[LoadQueue.scala 132:9:@13339.4]
  wire  storesToCheck_11_6; // @[LoadQueue.scala 131:10:@13340.4]
  wire  _T_10444; // @[LoadQueue.scala 131:81:@13343.4]
  wire  _T_10445; // @[LoadQueue.scala 131:72:@13344.4]
  wire  _T_10447; // @[LoadQueue.scala 132:33:@13345.4]
  wire  _T_10450; // @[LoadQueue.scala 132:41:@13347.4]
  wire  _T_10452; // @[LoadQueue.scala 132:9:@13348.4]
  wire  storesToCheck_11_7; // @[LoadQueue.scala 131:10:@13349.4]
  wire  _T_10458; // @[LoadQueue.scala 131:81:@13352.4]
  wire  _T_10459; // @[LoadQueue.scala 131:72:@13353.4]
  wire  _T_10461; // @[LoadQueue.scala 132:33:@13354.4]
  wire  _T_10464; // @[LoadQueue.scala 132:41:@13356.4]
  wire  _T_10466; // @[LoadQueue.scala 132:9:@13357.4]
  wire  storesToCheck_11_8; // @[LoadQueue.scala 131:10:@13358.4]
  wire  _T_10472; // @[LoadQueue.scala 131:81:@13361.4]
  wire  _T_10473; // @[LoadQueue.scala 131:72:@13362.4]
  wire  _T_10475; // @[LoadQueue.scala 132:33:@13363.4]
  wire  _T_10478; // @[LoadQueue.scala 132:41:@13365.4]
  wire  _T_10480; // @[LoadQueue.scala 132:9:@13366.4]
  wire  storesToCheck_11_9; // @[LoadQueue.scala 131:10:@13367.4]
  wire  _T_10486; // @[LoadQueue.scala 131:81:@13370.4]
  wire  _T_10487; // @[LoadQueue.scala 131:72:@13371.4]
  wire  _T_10489; // @[LoadQueue.scala 132:33:@13372.4]
  wire  _T_10492; // @[LoadQueue.scala 132:41:@13374.4]
  wire  _T_10494; // @[LoadQueue.scala 132:9:@13375.4]
  wire  storesToCheck_11_10; // @[LoadQueue.scala 131:10:@13376.4]
  wire  _T_10500; // @[LoadQueue.scala 131:81:@13379.4]
  wire  _T_10501; // @[LoadQueue.scala 131:72:@13380.4]
  wire  _T_10503; // @[LoadQueue.scala 132:33:@13381.4]
  wire  _T_10506; // @[LoadQueue.scala 132:41:@13383.4]
  wire  _T_10508; // @[LoadQueue.scala 132:9:@13384.4]
  wire  storesToCheck_11_11; // @[LoadQueue.scala 131:10:@13385.4]
  wire  _T_10514; // @[LoadQueue.scala 131:81:@13388.4]
  wire  _T_10515; // @[LoadQueue.scala 131:72:@13389.4]
  wire  _T_10517; // @[LoadQueue.scala 132:33:@13390.4]
  wire  _T_10520; // @[LoadQueue.scala 132:41:@13392.4]
  wire  _T_10522; // @[LoadQueue.scala 132:9:@13393.4]
  wire  storesToCheck_11_12; // @[LoadQueue.scala 131:10:@13394.4]
  wire  _T_10528; // @[LoadQueue.scala 131:81:@13397.4]
  wire  _T_10529; // @[LoadQueue.scala 131:72:@13398.4]
  wire  _T_10531; // @[LoadQueue.scala 132:33:@13399.4]
  wire  _T_10534; // @[LoadQueue.scala 132:41:@13401.4]
  wire  _T_10536; // @[LoadQueue.scala 132:9:@13402.4]
  wire  storesToCheck_11_13; // @[LoadQueue.scala 131:10:@13403.4]
  wire  _T_10542; // @[LoadQueue.scala 131:81:@13406.4]
  wire  _T_10543; // @[LoadQueue.scala 131:72:@13407.4]
  wire  _T_10545; // @[LoadQueue.scala 132:33:@13408.4]
  wire  _T_10548; // @[LoadQueue.scala 132:41:@13410.4]
  wire  _T_10550; // @[LoadQueue.scala 132:9:@13411.4]
  wire  storesToCheck_11_14; // @[LoadQueue.scala 131:10:@13412.4]
  wire  _T_10556; // @[LoadQueue.scala 131:81:@13415.4]
  wire  storesToCheck_11_15; // @[LoadQueue.scala 131:10:@13421.4]
  wire  storesToCheck_12_0; // @[LoadQueue.scala 131:10:@13463.4]
  wire  _T_10606; // @[LoadQueue.scala 131:81:@13466.4]
  wire  _T_10607; // @[LoadQueue.scala 131:72:@13467.4]
  wire  _T_10609; // @[LoadQueue.scala 132:33:@13468.4]
  wire  _T_10612; // @[LoadQueue.scala 132:41:@13470.4]
  wire  _T_10614; // @[LoadQueue.scala 132:9:@13471.4]
  wire  storesToCheck_12_1; // @[LoadQueue.scala 131:10:@13472.4]
  wire  _T_10620; // @[LoadQueue.scala 131:81:@13475.4]
  wire  _T_10621; // @[LoadQueue.scala 131:72:@13476.4]
  wire  _T_10623; // @[LoadQueue.scala 132:33:@13477.4]
  wire  _T_10626; // @[LoadQueue.scala 132:41:@13479.4]
  wire  _T_10628; // @[LoadQueue.scala 132:9:@13480.4]
  wire  storesToCheck_12_2; // @[LoadQueue.scala 131:10:@13481.4]
  wire  _T_10634; // @[LoadQueue.scala 131:81:@13484.4]
  wire  _T_10635; // @[LoadQueue.scala 131:72:@13485.4]
  wire  _T_10637; // @[LoadQueue.scala 132:33:@13486.4]
  wire  _T_10640; // @[LoadQueue.scala 132:41:@13488.4]
  wire  _T_10642; // @[LoadQueue.scala 132:9:@13489.4]
  wire  storesToCheck_12_3; // @[LoadQueue.scala 131:10:@13490.4]
  wire  _T_10648; // @[LoadQueue.scala 131:81:@13493.4]
  wire  _T_10649; // @[LoadQueue.scala 131:72:@13494.4]
  wire  _T_10651; // @[LoadQueue.scala 132:33:@13495.4]
  wire  _T_10654; // @[LoadQueue.scala 132:41:@13497.4]
  wire  _T_10656; // @[LoadQueue.scala 132:9:@13498.4]
  wire  storesToCheck_12_4; // @[LoadQueue.scala 131:10:@13499.4]
  wire  _T_10662; // @[LoadQueue.scala 131:81:@13502.4]
  wire  _T_10663; // @[LoadQueue.scala 131:72:@13503.4]
  wire  _T_10665; // @[LoadQueue.scala 132:33:@13504.4]
  wire  _T_10668; // @[LoadQueue.scala 132:41:@13506.4]
  wire  _T_10670; // @[LoadQueue.scala 132:9:@13507.4]
  wire  storesToCheck_12_5; // @[LoadQueue.scala 131:10:@13508.4]
  wire  _T_10676; // @[LoadQueue.scala 131:81:@13511.4]
  wire  _T_10677; // @[LoadQueue.scala 131:72:@13512.4]
  wire  _T_10679; // @[LoadQueue.scala 132:33:@13513.4]
  wire  _T_10682; // @[LoadQueue.scala 132:41:@13515.4]
  wire  _T_10684; // @[LoadQueue.scala 132:9:@13516.4]
  wire  storesToCheck_12_6; // @[LoadQueue.scala 131:10:@13517.4]
  wire  _T_10690; // @[LoadQueue.scala 131:81:@13520.4]
  wire  _T_10691; // @[LoadQueue.scala 131:72:@13521.4]
  wire  _T_10693; // @[LoadQueue.scala 132:33:@13522.4]
  wire  _T_10696; // @[LoadQueue.scala 132:41:@13524.4]
  wire  _T_10698; // @[LoadQueue.scala 132:9:@13525.4]
  wire  storesToCheck_12_7; // @[LoadQueue.scala 131:10:@13526.4]
  wire  _T_10704; // @[LoadQueue.scala 131:81:@13529.4]
  wire  _T_10705; // @[LoadQueue.scala 131:72:@13530.4]
  wire  _T_10707; // @[LoadQueue.scala 132:33:@13531.4]
  wire  _T_10710; // @[LoadQueue.scala 132:41:@13533.4]
  wire  _T_10712; // @[LoadQueue.scala 132:9:@13534.4]
  wire  storesToCheck_12_8; // @[LoadQueue.scala 131:10:@13535.4]
  wire  _T_10718; // @[LoadQueue.scala 131:81:@13538.4]
  wire  _T_10719; // @[LoadQueue.scala 131:72:@13539.4]
  wire  _T_10721; // @[LoadQueue.scala 132:33:@13540.4]
  wire  _T_10724; // @[LoadQueue.scala 132:41:@13542.4]
  wire  _T_10726; // @[LoadQueue.scala 132:9:@13543.4]
  wire  storesToCheck_12_9; // @[LoadQueue.scala 131:10:@13544.4]
  wire  _T_10732; // @[LoadQueue.scala 131:81:@13547.4]
  wire  _T_10733; // @[LoadQueue.scala 131:72:@13548.4]
  wire  _T_10735; // @[LoadQueue.scala 132:33:@13549.4]
  wire  _T_10738; // @[LoadQueue.scala 132:41:@13551.4]
  wire  _T_10740; // @[LoadQueue.scala 132:9:@13552.4]
  wire  storesToCheck_12_10; // @[LoadQueue.scala 131:10:@13553.4]
  wire  _T_10746; // @[LoadQueue.scala 131:81:@13556.4]
  wire  _T_10747; // @[LoadQueue.scala 131:72:@13557.4]
  wire  _T_10749; // @[LoadQueue.scala 132:33:@13558.4]
  wire  _T_10752; // @[LoadQueue.scala 132:41:@13560.4]
  wire  _T_10754; // @[LoadQueue.scala 132:9:@13561.4]
  wire  storesToCheck_12_11; // @[LoadQueue.scala 131:10:@13562.4]
  wire  _T_10760; // @[LoadQueue.scala 131:81:@13565.4]
  wire  _T_10761; // @[LoadQueue.scala 131:72:@13566.4]
  wire  _T_10763; // @[LoadQueue.scala 132:33:@13567.4]
  wire  _T_10766; // @[LoadQueue.scala 132:41:@13569.4]
  wire  _T_10768; // @[LoadQueue.scala 132:9:@13570.4]
  wire  storesToCheck_12_12; // @[LoadQueue.scala 131:10:@13571.4]
  wire  _T_10774; // @[LoadQueue.scala 131:81:@13574.4]
  wire  _T_10775; // @[LoadQueue.scala 131:72:@13575.4]
  wire  _T_10777; // @[LoadQueue.scala 132:33:@13576.4]
  wire  _T_10780; // @[LoadQueue.scala 132:41:@13578.4]
  wire  _T_10782; // @[LoadQueue.scala 132:9:@13579.4]
  wire  storesToCheck_12_13; // @[LoadQueue.scala 131:10:@13580.4]
  wire  _T_10788; // @[LoadQueue.scala 131:81:@13583.4]
  wire  _T_10789; // @[LoadQueue.scala 131:72:@13584.4]
  wire  _T_10791; // @[LoadQueue.scala 132:33:@13585.4]
  wire  _T_10794; // @[LoadQueue.scala 132:41:@13587.4]
  wire  _T_10796; // @[LoadQueue.scala 132:9:@13588.4]
  wire  storesToCheck_12_14; // @[LoadQueue.scala 131:10:@13589.4]
  wire  _T_10802; // @[LoadQueue.scala 131:81:@13592.4]
  wire  storesToCheck_12_15; // @[LoadQueue.scala 131:10:@13598.4]
  wire  storesToCheck_13_0; // @[LoadQueue.scala 131:10:@13640.4]
  wire  _T_10852; // @[LoadQueue.scala 131:81:@13643.4]
  wire  _T_10853; // @[LoadQueue.scala 131:72:@13644.4]
  wire  _T_10855; // @[LoadQueue.scala 132:33:@13645.4]
  wire  _T_10858; // @[LoadQueue.scala 132:41:@13647.4]
  wire  _T_10860; // @[LoadQueue.scala 132:9:@13648.4]
  wire  storesToCheck_13_1; // @[LoadQueue.scala 131:10:@13649.4]
  wire  _T_10866; // @[LoadQueue.scala 131:81:@13652.4]
  wire  _T_10867; // @[LoadQueue.scala 131:72:@13653.4]
  wire  _T_10869; // @[LoadQueue.scala 132:33:@13654.4]
  wire  _T_10872; // @[LoadQueue.scala 132:41:@13656.4]
  wire  _T_10874; // @[LoadQueue.scala 132:9:@13657.4]
  wire  storesToCheck_13_2; // @[LoadQueue.scala 131:10:@13658.4]
  wire  _T_10880; // @[LoadQueue.scala 131:81:@13661.4]
  wire  _T_10881; // @[LoadQueue.scala 131:72:@13662.4]
  wire  _T_10883; // @[LoadQueue.scala 132:33:@13663.4]
  wire  _T_10886; // @[LoadQueue.scala 132:41:@13665.4]
  wire  _T_10888; // @[LoadQueue.scala 132:9:@13666.4]
  wire  storesToCheck_13_3; // @[LoadQueue.scala 131:10:@13667.4]
  wire  _T_10894; // @[LoadQueue.scala 131:81:@13670.4]
  wire  _T_10895; // @[LoadQueue.scala 131:72:@13671.4]
  wire  _T_10897; // @[LoadQueue.scala 132:33:@13672.4]
  wire  _T_10900; // @[LoadQueue.scala 132:41:@13674.4]
  wire  _T_10902; // @[LoadQueue.scala 132:9:@13675.4]
  wire  storesToCheck_13_4; // @[LoadQueue.scala 131:10:@13676.4]
  wire  _T_10908; // @[LoadQueue.scala 131:81:@13679.4]
  wire  _T_10909; // @[LoadQueue.scala 131:72:@13680.4]
  wire  _T_10911; // @[LoadQueue.scala 132:33:@13681.4]
  wire  _T_10914; // @[LoadQueue.scala 132:41:@13683.4]
  wire  _T_10916; // @[LoadQueue.scala 132:9:@13684.4]
  wire  storesToCheck_13_5; // @[LoadQueue.scala 131:10:@13685.4]
  wire  _T_10922; // @[LoadQueue.scala 131:81:@13688.4]
  wire  _T_10923; // @[LoadQueue.scala 131:72:@13689.4]
  wire  _T_10925; // @[LoadQueue.scala 132:33:@13690.4]
  wire  _T_10928; // @[LoadQueue.scala 132:41:@13692.4]
  wire  _T_10930; // @[LoadQueue.scala 132:9:@13693.4]
  wire  storesToCheck_13_6; // @[LoadQueue.scala 131:10:@13694.4]
  wire  _T_10936; // @[LoadQueue.scala 131:81:@13697.4]
  wire  _T_10937; // @[LoadQueue.scala 131:72:@13698.4]
  wire  _T_10939; // @[LoadQueue.scala 132:33:@13699.4]
  wire  _T_10942; // @[LoadQueue.scala 132:41:@13701.4]
  wire  _T_10944; // @[LoadQueue.scala 132:9:@13702.4]
  wire  storesToCheck_13_7; // @[LoadQueue.scala 131:10:@13703.4]
  wire  _T_10950; // @[LoadQueue.scala 131:81:@13706.4]
  wire  _T_10951; // @[LoadQueue.scala 131:72:@13707.4]
  wire  _T_10953; // @[LoadQueue.scala 132:33:@13708.4]
  wire  _T_10956; // @[LoadQueue.scala 132:41:@13710.4]
  wire  _T_10958; // @[LoadQueue.scala 132:9:@13711.4]
  wire  storesToCheck_13_8; // @[LoadQueue.scala 131:10:@13712.4]
  wire  _T_10964; // @[LoadQueue.scala 131:81:@13715.4]
  wire  _T_10965; // @[LoadQueue.scala 131:72:@13716.4]
  wire  _T_10967; // @[LoadQueue.scala 132:33:@13717.4]
  wire  _T_10970; // @[LoadQueue.scala 132:41:@13719.4]
  wire  _T_10972; // @[LoadQueue.scala 132:9:@13720.4]
  wire  storesToCheck_13_9; // @[LoadQueue.scala 131:10:@13721.4]
  wire  _T_10978; // @[LoadQueue.scala 131:81:@13724.4]
  wire  _T_10979; // @[LoadQueue.scala 131:72:@13725.4]
  wire  _T_10981; // @[LoadQueue.scala 132:33:@13726.4]
  wire  _T_10984; // @[LoadQueue.scala 132:41:@13728.4]
  wire  _T_10986; // @[LoadQueue.scala 132:9:@13729.4]
  wire  storesToCheck_13_10; // @[LoadQueue.scala 131:10:@13730.4]
  wire  _T_10992; // @[LoadQueue.scala 131:81:@13733.4]
  wire  _T_10993; // @[LoadQueue.scala 131:72:@13734.4]
  wire  _T_10995; // @[LoadQueue.scala 132:33:@13735.4]
  wire  _T_10998; // @[LoadQueue.scala 132:41:@13737.4]
  wire  _T_11000; // @[LoadQueue.scala 132:9:@13738.4]
  wire  storesToCheck_13_11; // @[LoadQueue.scala 131:10:@13739.4]
  wire  _T_11006; // @[LoadQueue.scala 131:81:@13742.4]
  wire  _T_11007; // @[LoadQueue.scala 131:72:@13743.4]
  wire  _T_11009; // @[LoadQueue.scala 132:33:@13744.4]
  wire  _T_11012; // @[LoadQueue.scala 132:41:@13746.4]
  wire  _T_11014; // @[LoadQueue.scala 132:9:@13747.4]
  wire  storesToCheck_13_12; // @[LoadQueue.scala 131:10:@13748.4]
  wire  _T_11020; // @[LoadQueue.scala 131:81:@13751.4]
  wire  _T_11021; // @[LoadQueue.scala 131:72:@13752.4]
  wire  _T_11023; // @[LoadQueue.scala 132:33:@13753.4]
  wire  _T_11026; // @[LoadQueue.scala 132:41:@13755.4]
  wire  _T_11028; // @[LoadQueue.scala 132:9:@13756.4]
  wire  storesToCheck_13_13; // @[LoadQueue.scala 131:10:@13757.4]
  wire  _T_11034; // @[LoadQueue.scala 131:81:@13760.4]
  wire  _T_11035; // @[LoadQueue.scala 131:72:@13761.4]
  wire  _T_11037; // @[LoadQueue.scala 132:33:@13762.4]
  wire  _T_11040; // @[LoadQueue.scala 132:41:@13764.4]
  wire  _T_11042; // @[LoadQueue.scala 132:9:@13765.4]
  wire  storesToCheck_13_14; // @[LoadQueue.scala 131:10:@13766.4]
  wire  _T_11048; // @[LoadQueue.scala 131:81:@13769.4]
  wire  storesToCheck_13_15; // @[LoadQueue.scala 131:10:@13775.4]
  wire  storesToCheck_14_0; // @[LoadQueue.scala 131:10:@13817.4]
  wire  _T_11098; // @[LoadQueue.scala 131:81:@13820.4]
  wire  _T_11099; // @[LoadQueue.scala 131:72:@13821.4]
  wire  _T_11101; // @[LoadQueue.scala 132:33:@13822.4]
  wire  _T_11104; // @[LoadQueue.scala 132:41:@13824.4]
  wire  _T_11106; // @[LoadQueue.scala 132:9:@13825.4]
  wire  storesToCheck_14_1; // @[LoadQueue.scala 131:10:@13826.4]
  wire  _T_11112; // @[LoadQueue.scala 131:81:@13829.4]
  wire  _T_11113; // @[LoadQueue.scala 131:72:@13830.4]
  wire  _T_11115; // @[LoadQueue.scala 132:33:@13831.4]
  wire  _T_11118; // @[LoadQueue.scala 132:41:@13833.4]
  wire  _T_11120; // @[LoadQueue.scala 132:9:@13834.4]
  wire  storesToCheck_14_2; // @[LoadQueue.scala 131:10:@13835.4]
  wire  _T_11126; // @[LoadQueue.scala 131:81:@13838.4]
  wire  _T_11127; // @[LoadQueue.scala 131:72:@13839.4]
  wire  _T_11129; // @[LoadQueue.scala 132:33:@13840.4]
  wire  _T_11132; // @[LoadQueue.scala 132:41:@13842.4]
  wire  _T_11134; // @[LoadQueue.scala 132:9:@13843.4]
  wire  storesToCheck_14_3; // @[LoadQueue.scala 131:10:@13844.4]
  wire  _T_11140; // @[LoadQueue.scala 131:81:@13847.4]
  wire  _T_11141; // @[LoadQueue.scala 131:72:@13848.4]
  wire  _T_11143; // @[LoadQueue.scala 132:33:@13849.4]
  wire  _T_11146; // @[LoadQueue.scala 132:41:@13851.4]
  wire  _T_11148; // @[LoadQueue.scala 132:9:@13852.4]
  wire  storesToCheck_14_4; // @[LoadQueue.scala 131:10:@13853.4]
  wire  _T_11154; // @[LoadQueue.scala 131:81:@13856.4]
  wire  _T_11155; // @[LoadQueue.scala 131:72:@13857.4]
  wire  _T_11157; // @[LoadQueue.scala 132:33:@13858.4]
  wire  _T_11160; // @[LoadQueue.scala 132:41:@13860.4]
  wire  _T_11162; // @[LoadQueue.scala 132:9:@13861.4]
  wire  storesToCheck_14_5; // @[LoadQueue.scala 131:10:@13862.4]
  wire  _T_11168; // @[LoadQueue.scala 131:81:@13865.4]
  wire  _T_11169; // @[LoadQueue.scala 131:72:@13866.4]
  wire  _T_11171; // @[LoadQueue.scala 132:33:@13867.4]
  wire  _T_11174; // @[LoadQueue.scala 132:41:@13869.4]
  wire  _T_11176; // @[LoadQueue.scala 132:9:@13870.4]
  wire  storesToCheck_14_6; // @[LoadQueue.scala 131:10:@13871.4]
  wire  _T_11182; // @[LoadQueue.scala 131:81:@13874.4]
  wire  _T_11183; // @[LoadQueue.scala 131:72:@13875.4]
  wire  _T_11185; // @[LoadQueue.scala 132:33:@13876.4]
  wire  _T_11188; // @[LoadQueue.scala 132:41:@13878.4]
  wire  _T_11190; // @[LoadQueue.scala 132:9:@13879.4]
  wire  storesToCheck_14_7; // @[LoadQueue.scala 131:10:@13880.4]
  wire  _T_11196; // @[LoadQueue.scala 131:81:@13883.4]
  wire  _T_11197; // @[LoadQueue.scala 131:72:@13884.4]
  wire  _T_11199; // @[LoadQueue.scala 132:33:@13885.4]
  wire  _T_11202; // @[LoadQueue.scala 132:41:@13887.4]
  wire  _T_11204; // @[LoadQueue.scala 132:9:@13888.4]
  wire  storesToCheck_14_8; // @[LoadQueue.scala 131:10:@13889.4]
  wire  _T_11210; // @[LoadQueue.scala 131:81:@13892.4]
  wire  _T_11211; // @[LoadQueue.scala 131:72:@13893.4]
  wire  _T_11213; // @[LoadQueue.scala 132:33:@13894.4]
  wire  _T_11216; // @[LoadQueue.scala 132:41:@13896.4]
  wire  _T_11218; // @[LoadQueue.scala 132:9:@13897.4]
  wire  storesToCheck_14_9; // @[LoadQueue.scala 131:10:@13898.4]
  wire  _T_11224; // @[LoadQueue.scala 131:81:@13901.4]
  wire  _T_11225; // @[LoadQueue.scala 131:72:@13902.4]
  wire  _T_11227; // @[LoadQueue.scala 132:33:@13903.4]
  wire  _T_11230; // @[LoadQueue.scala 132:41:@13905.4]
  wire  _T_11232; // @[LoadQueue.scala 132:9:@13906.4]
  wire  storesToCheck_14_10; // @[LoadQueue.scala 131:10:@13907.4]
  wire  _T_11238; // @[LoadQueue.scala 131:81:@13910.4]
  wire  _T_11239; // @[LoadQueue.scala 131:72:@13911.4]
  wire  _T_11241; // @[LoadQueue.scala 132:33:@13912.4]
  wire  _T_11244; // @[LoadQueue.scala 132:41:@13914.4]
  wire  _T_11246; // @[LoadQueue.scala 132:9:@13915.4]
  wire  storesToCheck_14_11; // @[LoadQueue.scala 131:10:@13916.4]
  wire  _T_11252; // @[LoadQueue.scala 131:81:@13919.4]
  wire  _T_11253; // @[LoadQueue.scala 131:72:@13920.4]
  wire  _T_11255; // @[LoadQueue.scala 132:33:@13921.4]
  wire  _T_11258; // @[LoadQueue.scala 132:41:@13923.4]
  wire  _T_11260; // @[LoadQueue.scala 132:9:@13924.4]
  wire  storesToCheck_14_12; // @[LoadQueue.scala 131:10:@13925.4]
  wire  _T_11266; // @[LoadQueue.scala 131:81:@13928.4]
  wire  _T_11267; // @[LoadQueue.scala 131:72:@13929.4]
  wire  _T_11269; // @[LoadQueue.scala 132:33:@13930.4]
  wire  _T_11272; // @[LoadQueue.scala 132:41:@13932.4]
  wire  _T_11274; // @[LoadQueue.scala 132:9:@13933.4]
  wire  storesToCheck_14_13; // @[LoadQueue.scala 131:10:@13934.4]
  wire  _T_11280; // @[LoadQueue.scala 131:81:@13937.4]
  wire  _T_11281; // @[LoadQueue.scala 131:72:@13938.4]
  wire  _T_11283; // @[LoadQueue.scala 132:33:@13939.4]
  wire  _T_11286; // @[LoadQueue.scala 132:41:@13941.4]
  wire  _T_11288; // @[LoadQueue.scala 132:9:@13942.4]
  wire  storesToCheck_14_14; // @[LoadQueue.scala 131:10:@13943.4]
  wire  _T_11294; // @[LoadQueue.scala 131:81:@13946.4]
  wire  storesToCheck_14_15; // @[LoadQueue.scala 131:10:@13952.4]
  wire  storesToCheck_15_0; // @[LoadQueue.scala 131:10:@13994.4]
  wire  _T_11344; // @[LoadQueue.scala 131:81:@13997.4]
  wire  _T_11345; // @[LoadQueue.scala 131:72:@13998.4]
  wire  _T_11347; // @[LoadQueue.scala 132:33:@13999.4]
  wire  _T_11350; // @[LoadQueue.scala 132:41:@14001.4]
  wire  _T_11352; // @[LoadQueue.scala 132:9:@14002.4]
  wire  storesToCheck_15_1; // @[LoadQueue.scala 131:10:@14003.4]
  wire  _T_11358; // @[LoadQueue.scala 131:81:@14006.4]
  wire  _T_11359; // @[LoadQueue.scala 131:72:@14007.4]
  wire  _T_11361; // @[LoadQueue.scala 132:33:@14008.4]
  wire  _T_11364; // @[LoadQueue.scala 132:41:@14010.4]
  wire  _T_11366; // @[LoadQueue.scala 132:9:@14011.4]
  wire  storesToCheck_15_2; // @[LoadQueue.scala 131:10:@14012.4]
  wire  _T_11372; // @[LoadQueue.scala 131:81:@14015.4]
  wire  _T_11373; // @[LoadQueue.scala 131:72:@14016.4]
  wire  _T_11375; // @[LoadQueue.scala 132:33:@14017.4]
  wire  _T_11378; // @[LoadQueue.scala 132:41:@14019.4]
  wire  _T_11380; // @[LoadQueue.scala 132:9:@14020.4]
  wire  storesToCheck_15_3; // @[LoadQueue.scala 131:10:@14021.4]
  wire  _T_11386; // @[LoadQueue.scala 131:81:@14024.4]
  wire  _T_11387; // @[LoadQueue.scala 131:72:@14025.4]
  wire  _T_11389; // @[LoadQueue.scala 132:33:@14026.4]
  wire  _T_11392; // @[LoadQueue.scala 132:41:@14028.4]
  wire  _T_11394; // @[LoadQueue.scala 132:9:@14029.4]
  wire  storesToCheck_15_4; // @[LoadQueue.scala 131:10:@14030.4]
  wire  _T_11400; // @[LoadQueue.scala 131:81:@14033.4]
  wire  _T_11401; // @[LoadQueue.scala 131:72:@14034.4]
  wire  _T_11403; // @[LoadQueue.scala 132:33:@14035.4]
  wire  _T_11406; // @[LoadQueue.scala 132:41:@14037.4]
  wire  _T_11408; // @[LoadQueue.scala 132:9:@14038.4]
  wire  storesToCheck_15_5; // @[LoadQueue.scala 131:10:@14039.4]
  wire  _T_11414; // @[LoadQueue.scala 131:81:@14042.4]
  wire  _T_11415; // @[LoadQueue.scala 131:72:@14043.4]
  wire  _T_11417; // @[LoadQueue.scala 132:33:@14044.4]
  wire  _T_11420; // @[LoadQueue.scala 132:41:@14046.4]
  wire  _T_11422; // @[LoadQueue.scala 132:9:@14047.4]
  wire  storesToCheck_15_6; // @[LoadQueue.scala 131:10:@14048.4]
  wire  _T_11428; // @[LoadQueue.scala 131:81:@14051.4]
  wire  _T_11429; // @[LoadQueue.scala 131:72:@14052.4]
  wire  _T_11431; // @[LoadQueue.scala 132:33:@14053.4]
  wire  _T_11434; // @[LoadQueue.scala 132:41:@14055.4]
  wire  _T_11436; // @[LoadQueue.scala 132:9:@14056.4]
  wire  storesToCheck_15_7; // @[LoadQueue.scala 131:10:@14057.4]
  wire  _T_11442; // @[LoadQueue.scala 131:81:@14060.4]
  wire  _T_11443; // @[LoadQueue.scala 131:72:@14061.4]
  wire  _T_11445; // @[LoadQueue.scala 132:33:@14062.4]
  wire  _T_11448; // @[LoadQueue.scala 132:41:@14064.4]
  wire  _T_11450; // @[LoadQueue.scala 132:9:@14065.4]
  wire  storesToCheck_15_8; // @[LoadQueue.scala 131:10:@14066.4]
  wire  _T_11456; // @[LoadQueue.scala 131:81:@14069.4]
  wire  _T_11457; // @[LoadQueue.scala 131:72:@14070.4]
  wire  _T_11459; // @[LoadQueue.scala 132:33:@14071.4]
  wire  _T_11462; // @[LoadQueue.scala 132:41:@14073.4]
  wire  _T_11464; // @[LoadQueue.scala 132:9:@14074.4]
  wire  storesToCheck_15_9; // @[LoadQueue.scala 131:10:@14075.4]
  wire  _T_11470; // @[LoadQueue.scala 131:81:@14078.4]
  wire  _T_11471; // @[LoadQueue.scala 131:72:@14079.4]
  wire  _T_11473; // @[LoadQueue.scala 132:33:@14080.4]
  wire  _T_11476; // @[LoadQueue.scala 132:41:@14082.4]
  wire  _T_11478; // @[LoadQueue.scala 132:9:@14083.4]
  wire  storesToCheck_15_10; // @[LoadQueue.scala 131:10:@14084.4]
  wire  _T_11484; // @[LoadQueue.scala 131:81:@14087.4]
  wire  _T_11485; // @[LoadQueue.scala 131:72:@14088.4]
  wire  _T_11487; // @[LoadQueue.scala 132:33:@14089.4]
  wire  _T_11490; // @[LoadQueue.scala 132:41:@14091.4]
  wire  _T_11492; // @[LoadQueue.scala 132:9:@14092.4]
  wire  storesToCheck_15_11; // @[LoadQueue.scala 131:10:@14093.4]
  wire  _T_11498; // @[LoadQueue.scala 131:81:@14096.4]
  wire  _T_11499; // @[LoadQueue.scala 131:72:@14097.4]
  wire  _T_11501; // @[LoadQueue.scala 132:33:@14098.4]
  wire  _T_11504; // @[LoadQueue.scala 132:41:@14100.4]
  wire  _T_11506; // @[LoadQueue.scala 132:9:@14101.4]
  wire  storesToCheck_15_12; // @[LoadQueue.scala 131:10:@14102.4]
  wire  _T_11512; // @[LoadQueue.scala 131:81:@14105.4]
  wire  _T_11513; // @[LoadQueue.scala 131:72:@14106.4]
  wire  _T_11515; // @[LoadQueue.scala 132:33:@14107.4]
  wire  _T_11518; // @[LoadQueue.scala 132:41:@14109.4]
  wire  _T_11520; // @[LoadQueue.scala 132:9:@14110.4]
  wire  storesToCheck_15_13; // @[LoadQueue.scala 131:10:@14111.4]
  wire  _T_11526; // @[LoadQueue.scala 131:81:@14114.4]
  wire  _T_11527; // @[LoadQueue.scala 131:72:@14115.4]
  wire  _T_11529; // @[LoadQueue.scala 132:33:@14116.4]
  wire  _T_11532; // @[LoadQueue.scala 132:41:@14118.4]
  wire  _T_11534; // @[LoadQueue.scala 132:9:@14119.4]
  wire  storesToCheck_15_14; // @[LoadQueue.scala 131:10:@14120.4]
  wire  _T_11540; // @[LoadQueue.scala 131:81:@14123.4]
  wire  storesToCheck_15_15; // @[LoadQueue.scala 131:10:@14129.4]
  wire  _T_12802; // @[LoadQueue.scala 141:18:@14164.4]
  wire  entriesToCheck_0_0; // @[LoadQueue.scala 141:26:@14165.4]
  wire  _T_12804; // @[LoadQueue.scala 141:18:@14166.4]
  wire  entriesToCheck_0_1; // @[LoadQueue.scala 141:26:@14167.4]
  wire  _T_12806; // @[LoadQueue.scala 141:18:@14168.4]
  wire  entriesToCheck_0_2; // @[LoadQueue.scala 141:26:@14169.4]
  wire  _T_12808; // @[LoadQueue.scala 141:18:@14170.4]
  wire  entriesToCheck_0_3; // @[LoadQueue.scala 141:26:@14171.4]
  wire  _T_12810; // @[LoadQueue.scala 141:18:@14172.4]
  wire  entriesToCheck_0_4; // @[LoadQueue.scala 141:26:@14173.4]
  wire  _T_12812; // @[LoadQueue.scala 141:18:@14174.4]
  wire  entriesToCheck_0_5; // @[LoadQueue.scala 141:26:@14175.4]
  wire  _T_12814; // @[LoadQueue.scala 141:18:@14176.4]
  wire  entriesToCheck_0_6; // @[LoadQueue.scala 141:26:@14177.4]
  wire  _T_12816; // @[LoadQueue.scala 141:18:@14178.4]
  wire  entriesToCheck_0_7; // @[LoadQueue.scala 141:26:@14179.4]
  wire  _T_12818; // @[LoadQueue.scala 141:18:@14180.4]
  wire  entriesToCheck_0_8; // @[LoadQueue.scala 141:26:@14181.4]
  wire  _T_12820; // @[LoadQueue.scala 141:18:@14182.4]
  wire  entriesToCheck_0_9; // @[LoadQueue.scala 141:26:@14183.4]
  wire  _T_12822; // @[LoadQueue.scala 141:18:@14184.4]
  wire  entriesToCheck_0_10; // @[LoadQueue.scala 141:26:@14185.4]
  wire  _T_12824; // @[LoadQueue.scala 141:18:@14186.4]
  wire  entriesToCheck_0_11; // @[LoadQueue.scala 141:26:@14187.4]
  wire  _T_12826; // @[LoadQueue.scala 141:18:@14188.4]
  wire  entriesToCheck_0_12; // @[LoadQueue.scala 141:26:@14189.4]
  wire  _T_12828; // @[LoadQueue.scala 141:18:@14190.4]
  wire  entriesToCheck_0_13; // @[LoadQueue.scala 141:26:@14191.4]
  wire  _T_12830; // @[LoadQueue.scala 141:18:@14192.4]
  wire  entriesToCheck_0_14; // @[LoadQueue.scala 141:26:@14193.4]
  wire  _T_12832; // @[LoadQueue.scala 141:18:@14194.4]
  wire  entriesToCheck_0_15; // @[LoadQueue.scala 141:26:@14195.4]
  wire  _T_12834; // @[LoadQueue.scala 141:18:@14212.4]
  wire  entriesToCheck_1_0; // @[LoadQueue.scala 141:26:@14213.4]
  wire  _T_12836; // @[LoadQueue.scala 141:18:@14214.4]
  wire  entriesToCheck_1_1; // @[LoadQueue.scala 141:26:@14215.4]
  wire  _T_12838; // @[LoadQueue.scala 141:18:@14216.4]
  wire  entriesToCheck_1_2; // @[LoadQueue.scala 141:26:@14217.4]
  wire  _T_12840; // @[LoadQueue.scala 141:18:@14218.4]
  wire  entriesToCheck_1_3; // @[LoadQueue.scala 141:26:@14219.4]
  wire  _T_12842; // @[LoadQueue.scala 141:18:@14220.4]
  wire  entriesToCheck_1_4; // @[LoadQueue.scala 141:26:@14221.4]
  wire  _T_12844; // @[LoadQueue.scala 141:18:@14222.4]
  wire  entriesToCheck_1_5; // @[LoadQueue.scala 141:26:@14223.4]
  wire  _T_12846; // @[LoadQueue.scala 141:18:@14224.4]
  wire  entriesToCheck_1_6; // @[LoadQueue.scala 141:26:@14225.4]
  wire  _T_12848; // @[LoadQueue.scala 141:18:@14226.4]
  wire  entriesToCheck_1_7; // @[LoadQueue.scala 141:26:@14227.4]
  wire  _T_12850; // @[LoadQueue.scala 141:18:@14228.4]
  wire  entriesToCheck_1_8; // @[LoadQueue.scala 141:26:@14229.4]
  wire  _T_12852; // @[LoadQueue.scala 141:18:@14230.4]
  wire  entriesToCheck_1_9; // @[LoadQueue.scala 141:26:@14231.4]
  wire  _T_12854; // @[LoadQueue.scala 141:18:@14232.4]
  wire  entriesToCheck_1_10; // @[LoadQueue.scala 141:26:@14233.4]
  wire  _T_12856; // @[LoadQueue.scala 141:18:@14234.4]
  wire  entriesToCheck_1_11; // @[LoadQueue.scala 141:26:@14235.4]
  wire  _T_12858; // @[LoadQueue.scala 141:18:@14236.4]
  wire  entriesToCheck_1_12; // @[LoadQueue.scala 141:26:@14237.4]
  wire  _T_12860; // @[LoadQueue.scala 141:18:@14238.4]
  wire  entriesToCheck_1_13; // @[LoadQueue.scala 141:26:@14239.4]
  wire  _T_12862; // @[LoadQueue.scala 141:18:@14240.4]
  wire  entriesToCheck_1_14; // @[LoadQueue.scala 141:26:@14241.4]
  wire  _T_12864; // @[LoadQueue.scala 141:18:@14242.4]
  wire  entriesToCheck_1_15; // @[LoadQueue.scala 141:26:@14243.4]
  wire  _T_12866; // @[LoadQueue.scala 141:18:@14260.4]
  wire  entriesToCheck_2_0; // @[LoadQueue.scala 141:26:@14261.4]
  wire  _T_12868; // @[LoadQueue.scala 141:18:@14262.4]
  wire  entriesToCheck_2_1; // @[LoadQueue.scala 141:26:@14263.4]
  wire  _T_12870; // @[LoadQueue.scala 141:18:@14264.4]
  wire  entriesToCheck_2_2; // @[LoadQueue.scala 141:26:@14265.4]
  wire  _T_12872; // @[LoadQueue.scala 141:18:@14266.4]
  wire  entriesToCheck_2_3; // @[LoadQueue.scala 141:26:@14267.4]
  wire  _T_12874; // @[LoadQueue.scala 141:18:@14268.4]
  wire  entriesToCheck_2_4; // @[LoadQueue.scala 141:26:@14269.4]
  wire  _T_12876; // @[LoadQueue.scala 141:18:@14270.4]
  wire  entriesToCheck_2_5; // @[LoadQueue.scala 141:26:@14271.4]
  wire  _T_12878; // @[LoadQueue.scala 141:18:@14272.4]
  wire  entriesToCheck_2_6; // @[LoadQueue.scala 141:26:@14273.4]
  wire  _T_12880; // @[LoadQueue.scala 141:18:@14274.4]
  wire  entriesToCheck_2_7; // @[LoadQueue.scala 141:26:@14275.4]
  wire  _T_12882; // @[LoadQueue.scala 141:18:@14276.4]
  wire  entriesToCheck_2_8; // @[LoadQueue.scala 141:26:@14277.4]
  wire  _T_12884; // @[LoadQueue.scala 141:18:@14278.4]
  wire  entriesToCheck_2_9; // @[LoadQueue.scala 141:26:@14279.4]
  wire  _T_12886; // @[LoadQueue.scala 141:18:@14280.4]
  wire  entriesToCheck_2_10; // @[LoadQueue.scala 141:26:@14281.4]
  wire  _T_12888; // @[LoadQueue.scala 141:18:@14282.4]
  wire  entriesToCheck_2_11; // @[LoadQueue.scala 141:26:@14283.4]
  wire  _T_12890; // @[LoadQueue.scala 141:18:@14284.4]
  wire  entriesToCheck_2_12; // @[LoadQueue.scala 141:26:@14285.4]
  wire  _T_12892; // @[LoadQueue.scala 141:18:@14286.4]
  wire  entriesToCheck_2_13; // @[LoadQueue.scala 141:26:@14287.4]
  wire  _T_12894; // @[LoadQueue.scala 141:18:@14288.4]
  wire  entriesToCheck_2_14; // @[LoadQueue.scala 141:26:@14289.4]
  wire  _T_12896; // @[LoadQueue.scala 141:18:@14290.4]
  wire  entriesToCheck_2_15; // @[LoadQueue.scala 141:26:@14291.4]
  wire  _T_12898; // @[LoadQueue.scala 141:18:@14308.4]
  wire  entriesToCheck_3_0; // @[LoadQueue.scala 141:26:@14309.4]
  wire  _T_12900; // @[LoadQueue.scala 141:18:@14310.4]
  wire  entriesToCheck_3_1; // @[LoadQueue.scala 141:26:@14311.4]
  wire  _T_12902; // @[LoadQueue.scala 141:18:@14312.4]
  wire  entriesToCheck_3_2; // @[LoadQueue.scala 141:26:@14313.4]
  wire  _T_12904; // @[LoadQueue.scala 141:18:@14314.4]
  wire  entriesToCheck_3_3; // @[LoadQueue.scala 141:26:@14315.4]
  wire  _T_12906; // @[LoadQueue.scala 141:18:@14316.4]
  wire  entriesToCheck_3_4; // @[LoadQueue.scala 141:26:@14317.4]
  wire  _T_12908; // @[LoadQueue.scala 141:18:@14318.4]
  wire  entriesToCheck_3_5; // @[LoadQueue.scala 141:26:@14319.4]
  wire  _T_12910; // @[LoadQueue.scala 141:18:@14320.4]
  wire  entriesToCheck_3_6; // @[LoadQueue.scala 141:26:@14321.4]
  wire  _T_12912; // @[LoadQueue.scala 141:18:@14322.4]
  wire  entriesToCheck_3_7; // @[LoadQueue.scala 141:26:@14323.4]
  wire  _T_12914; // @[LoadQueue.scala 141:18:@14324.4]
  wire  entriesToCheck_3_8; // @[LoadQueue.scala 141:26:@14325.4]
  wire  _T_12916; // @[LoadQueue.scala 141:18:@14326.4]
  wire  entriesToCheck_3_9; // @[LoadQueue.scala 141:26:@14327.4]
  wire  _T_12918; // @[LoadQueue.scala 141:18:@14328.4]
  wire  entriesToCheck_3_10; // @[LoadQueue.scala 141:26:@14329.4]
  wire  _T_12920; // @[LoadQueue.scala 141:18:@14330.4]
  wire  entriesToCheck_3_11; // @[LoadQueue.scala 141:26:@14331.4]
  wire  _T_12922; // @[LoadQueue.scala 141:18:@14332.4]
  wire  entriesToCheck_3_12; // @[LoadQueue.scala 141:26:@14333.4]
  wire  _T_12924; // @[LoadQueue.scala 141:18:@14334.4]
  wire  entriesToCheck_3_13; // @[LoadQueue.scala 141:26:@14335.4]
  wire  _T_12926; // @[LoadQueue.scala 141:18:@14336.4]
  wire  entriesToCheck_3_14; // @[LoadQueue.scala 141:26:@14337.4]
  wire  _T_12928; // @[LoadQueue.scala 141:18:@14338.4]
  wire  entriesToCheck_3_15; // @[LoadQueue.scala 141:26:@14339.4]
  wire  _T_12930; // @[LoadQueue.scala 141:18:@14356.4]
  wire  entriesToCheck_4_0; // @[LoadQueue.scala 141:26:@14357.4]
  wire  _T_12932; // @[LoadQueue.scala 141:18:@14358.4]
  wire  entriesToCheck_4_1; // @[LoadQueue.scala 141:26:@14359.4]
  wire  _T_12934; // @[LoadQueue.scala 141:18:@14360.4]
  wire  entriesToCheck_4_2; // @[LoadQueue.scala 141:26:@14361.4]
  wire  _T_12936; // @[LoadQueue.scala 141:18:@14362.4]
  wire  entriesToCheck_4_3; // @[LoadQueue.scala 141:26:@14363.4]
  wire  _T_12938; // @[LoadQueue.scala 141:18:@14364.4]
  wire  entriesToCheck_4_4; // @[LoadQueue.scala 141:26:@14365.4]
  wire  _T_12940; // @[LoadQueue.scala 141:18:@14366.4]
  wire  entriesToCheck_4_5; // @[LoadQueue.scala 141:26:@14367.4]
  wire  _T_12942; // @[LoadQueue.scala 141:18:@14368.4]
  wire  entriesToCheck_4_6; // @[LoadQueue.scala 141:26:@14369.4]
  wire  _T_12944; // @[LoadQueue.scala 141:18:@14370.4]
  wire  entriesToCheck_4_7; // @[LoadQueue.scala 141:26:@14371.4]
  wire  _T_12946; // @[LoadQueue.scala 141:18:@14372.4]
  wire  entriesToCheck_4_8; // @[LoadQueue.scala 141:26:@14373.4]
  wire  _T_12948; // @[LoadQueue.scala 141:18:@14374.4]
  wire  entriesToCheck_4_9; // @[LoadQueue.scala 141:26:@14375.4]
  wire  _T_12950; // @[LoadQueue.scala 141:18:@14376.4]
  wire  entriesToCheck_4_10; // @[LoadQueue.scala 141:26:@14377.4]
  wire  _T_12952; // @[LoadQueue.scala 141:18:@14378.4]
  wire  entriesToCheck_4_11; // @[LoadQueue.scala 141:26:@14379.4]
  wire  _T_12954; // @[LoadQueue.scala 141:18:@14380.4]
  wire  entriesToCheck_4_12; // @[LoadQueue.scala 141:26:@14381.4]
  wire  _T_12956; // @[LoadQueue.scala 141:18:@14382.4]
  wire  entriesToCheck_4_13; // @[LoadQueue.scala 141:26:@14383.4]
  wire  _T_12958; // @[LoadQueue.scala 141:18:@14384.4]
  wire  entriesToCheck_4_14; // @[LoadQueue.scala 141:26:@14385.4]
  wire  _T_12960; // @[LoadQueue.scala 141:18:@14386.4]
  wire  entriesToCheck_4_15; // @[LoadQueue.scala 141:26:@14387.4]
  wire  _T_12962; // @[LoadQueue.scala 141:18:@14404.4]
  wire  entriesToCheck_5_0; // @[LoadQueue.scala 141:26:@14405.4]
  wire  _T_12964; // @[LoadQueue.scala 141:18:@14406.4]
  wire  entriesToCheck_5_1; // @[LoadQueue.scala 141:26:@14407.4]
  wire  _T_12966; // @[LoadQueue.scala 141:18:@14408.4]
  wire  entriesToCheck_5_2; // @[LoadQueue.scala 141:26:@14409.4]
  wire  _T_12968; // @[LoadQueue.scala 141:18:@14410.4]
  wire  entriesToCheck_5_3; // @[LoadQueue.scala 141:26:@14411.4]
  wire  _T_12970; // @[LoadQueue.scala 141:18:@14412.4]
  wire  entriesToCheck_5_4; // @[LoadQueue.scala 141:26:@14413.4]
  wire  _T_12972; // @[LoadQueue.scala 141:18:@14414.4]
  wire  entriesToCheck_5_5; // @[LoadQueue.scala 141:26:@14415.4]
  wire  _T_12974; // @[LoadQueue.scala 141:18:@14416.4]
  wire  entriesToCheck_5_6; // @[LoadQueue.scala 141:26:@14417.4]
  wire  _T_12976; // @[LoadQueue.scala 141:18:@14418.4]
  wire  entriesToCheck_5_7; // @[LoadQueue.scala 141:26:@14419.4]
  wire  _T_12978; // @[LoadQueue.scala 141:18:@14420.4]
  wire  entriesToCheck_5_8; // @[LoadQueue.scala 141:26:@14421.4]
  wire  _T_12980; // @[LoadQueue.scala 141:18:@14422.4]
  wire  entriesToCheck_5_9; // @[LoadQueue.scala 141:26:@14423.4]
  wire  _T_12982; // @[LoadQueue.scala 141:18:@14424.4]
  wire  entriesToCheck_5_10; // @[LoadQueue.scala 141:26:@14425.4]
  wire  _T_12984; // @[LoadQueue.scala 141:18:@14426.4]
  wire  entriesToCheck_5_11; // @[LoadQueue.scala 141:26:@14427.4]
  wire  _T_12986; // @[LoadQueue.scala 141:18:@14428.4]
  wire  entriesToCheck_5_12; // @[LoadQueue.scala 141:26:@14429.4]
  wire  _T_12988; // @[LoadQueue.scala 141:18:@14430.4]
  wire  entriesToCheck_5_13; // @[LoadQueue.scala 141:26:@14431.4]
  wire  _T_12990; // @[LoadQueue.scala 141:18:@14432.4]
  wire  entriesToCheck_5_14; // @[LoadQueue.scala 141:26:@14433.4]
  wire  _T_12992; // @[LoadQueue.scala 141:18:@14434.4]
  wire  entriesToCheck_5_15; // @[LoadQueue.scala 141:26:@14435.4]
  wire  _T_12994; // @[LoadQueue.scala 141:18:@14452.4]
  wire  entriesToCheck_6_0; // @[LoadQueue.scala 141:26:@14453.4]
  wire  _T_12996; // @[LoadQueue.scala 141:18:@14454.4]
  wire  entriesToCheck_6_1; // @[LoadQueue.scala 141:26:@14455.4]
  wire  _T_12998; // @[LoadQueue.scala 141:18:@14456.4]
  wire  entriesToCheck_6_2; // @[LoadQueue.scala 141:26:@14457.4]
  wire  _T_13000; // @[LoadQueue.scala 141:18:@14458.4]
  wire  entriesToCheck_6_3; // @[LoadQueue.scala 141:26:@14459.4]
  wire  _T_13002; // @[LoadQueue.scala 141:18:@14460.4]
  wire  entriesToCheck_6_4; // @[LoadQueue.scala 141:26:@14461.4]
  wire  _T_13004; // @[LoadQueue.scala 141:18:@14462.4]
  wire  entriesToCheck_6_5; // @[LoadQueue.scala 141:26:@14463.4]
  wire  _T_13006; // @[LoadQueue.scala 141:18:@14464.4]
  wire  entriesToCheck_6_6; // @[LoadQueue.scala 141:26:@14465.4]
  wire  _T_13008; // @[LoadQueue.scala 141:18:@14466.4]
  wire  entriesToCheck_6_7; // @[LoadQueue.scala 141:26:@14467.4]
  wire  _T_13010; // @[LoadQueue.scala 141:18:@14468.4]
  wire  entriesToCheck_6_8; // @[LoadQueue.scala 141:26:@14469.4]
  wire  _T_13012; // @[LoadQueue.scala 141:18:@14470.4]
  wire  entriesToCheck_6_9; // @[LoadQueue.scala 141:26:@14471.4]
  wire  _T_13014; // @[LoadQueue.scala 141:18:@14472.4]
  wire  entriesToCheck_6_10; // @[LoadQueue.scala 141:26:@14473.4]
  wire  _T_13016; // @[LoadQueue.scala 141:18:@14474.4]
  wire  entriesToCheck_6_11; // @[LoadQueue.scala 141:26:@14475.4]
  wire  _T_13018; // @[LoadQueue.scala 141:18:@14476.4]
  wire  entriesToCheck_6_12; // @[LoadQueue.scala 141:26:@14477.4]
  wire  _T_13020; // @[LoadQueue.scala 141:18:@14478.4]
  wire  entriesToCheck_6_13; // @[LoadQueue.scala 141:26:@14479.4]
  wire  _T_13022; // @[LoadQueue.scala 141:18:@14480.4]
  wire  entriesToCheck_6_14; // @[LoadQueue.scala 141:26:@14481.4]
  wire  _T_13024; // @[LoadQueue.scala 141:18:@14482.4]
  wire  entriesToCheck_6_15; // @[LoadQueue.scala 141:26:@14483.4]
  wire  _T_13026; // @[LoadQueue.scala 141:18:@14500.4]
  wire  entriesToCheck_7_0; // @[LoadQueue.scala 141:26:@14501.4]
  wire  _T_13028; // @[LoadQueue.scala 141:18:@14502.4]
  wire  entriesToCheck_7_1; // @[LoadQueue.scala 141:26:@14503.4]
  wire  _T_13030; // @[LoadQueue.scala 141:18:@14504.4]
  wire  entriesToCheck_7_2; // @[LoadQueue.scala 141:26:@14505.4]
  wire  _T_13032; // @[LoadQueue.scala 141:18:@14506.4]
  wire  entriesToCheck_7_3; // @[LoadQueue.scala 141:26:@14507.4]
  wire  _T_13034; // @[LoadQueue.scala 141:18:@14508.4]
  wire  entriesToCheck_7_4; // @[LoadQueue.scala 141:26:@14509.4]
  wire  _T_13036; // @[LoadQueue.scala 141:18:@14510.4]
  wire  entriesToCheck_7_5; // @[LoadQueue.scala 141:26:@14511.4]
  wire  _T_13038; // @[LoadQueue.scala 141:18:@14512.4]
  wire  entriesToCheck_7_6; // @[LoadQueue.scala 141:26:@14513.4]
  wire  _T_13040; // @[LoadQueue.scala 141:18:@14514.4]
  wire  entriesToCheck_7_7; // @[LoadQueue.scala 141:26:@14515.4]
  wire  _T_13042; // @[LoadQueue.scala 141:18:@14516.4]
  wire  entriesToCheck_7_8; // @[LoadQueue.scala 141:26:@14517.4]
  wire  _T_13044; // @[LoadQueue.scala 141:18:@14518.4]
  wire  entriesToCheck_7_9; // @[LoadQueue.scala 141:26:@14519.4]
  wire  _T_13046; // @[LoadQueue.scala 141:18:@14520.4]
  wire  entriesToCheck_7_10; // @[LoadQueue.scala 141:26:@14521.4]
  wire  _T_13048; // @[LoadQueue.scala 141:18:@14522.4]
  wire  entriesToCheck_7_11; // @[LoadQueue.scala 141:26:@14523.4]
  wire  _T_13050; // @[LoadQueue.scala 141:18:@14524.4]
  wire  entriesToCheck_7_12; // @[LoadQueue.scala 141:26:@14525.4]
  wire  _T_13052; // @[LoadQueue.scala 141:18:@14526.4]
  wire  entriesToCheck_7_13; // @[LoadQueue.scala 141:26:@14527.4]
  wire  _T_13054; // @[LoadQueue.scala 141:18:@14528.4]
  wire  entriesToCheck_7_14; // @[LoadQueue.scala 141:26:@14529.4]
  wire  _T_13056; // @[LoadQueue.scala 141:18:@14530.4]
  wire  entriesToCheck_7_15; // @[LoadQueue.scala 141:26:@14531.4]
  wire  _T_13058; // @[LoadQueue.scala 141:18:@14548.4]
  wire  entriesToCheck_8_0; // @[LoadQueue.scala 141:26:@14549.4]
  wire  _T_13060; // @[LoadQueue.scala 141:18:@14550.4]
  wire  entriesToCheck_8_1; // @[LoadQueue.scala 141:26:@14551.4]
  wire  _T_13062; // @[LoadQueue.scala 141:18:@14552.4]
  wire  entriesToCheck_8_2; // @[LoadQueue.scala 141:26:@14553.4]
  wire  _T_13064; // @[LoadQueue.scala 141:18:@14554.4]
  wire  entriesToCheck_8_3; // @[LoadQueue.scala 141:26:@14555.4]
  wire  _T_13066; // @[LoadQueue.scala 141:18:@14556.4]
  wire  entriesToCheck_8_4; // @[LoadQueue.scala 141:26:@14557.4]
  wire  _T_13068; // @[LoadQueue.scala 141:18:@14558.4]
  wire  entriesToCheck_8_5; // @[LoadQueue.scala 141:26:@14559.4]
  wire  _T_13070; // @[LoadQueue.scala 141:18:@14560.4]
  wire  entriesToCheck_8_6; // @[LoadQueue.scala 141:26:@14561.4]
  wire  _T_13072; // @[LoadQueue.scala 141:18:@14562.4]
  wire  entriesToCheck_8_7; // @[LoadQueue.scala 141:26:@14563.4]
  wire  _T_13074; // @[LoadQueue.scala 141:18:@14564.4]
  wire  entriesToCheck_8_8; // @[LoadQueue.scala 141:26:@14565.4]
  wire  _T_13076; // @[LoadQueue.scala 141:18:@14566.4]
  wire  entriesToCheck_8_9; // @[LoadQueue.scala 141:26:@14567.4]
  wire  _T_13078; // @[LoadQueue.scala 141:18:@14568.4]
  wire  entriesToCheck_8_10; // @[LoadQueue.scala 141:26:@14569.4]
  wire  _T_13080; // @[LoadQueue.scala 141:18:@14570.4]
  wire  entriesToCheck_8_11; // @[LoadQueue.scala 141:26:@14571.4]
  wire  _T_13082; // @[LoadQueue.scala 141:18:@14572.4]
  wire  entriesToCheck_8_12; // @[LoadQueue.scala 141:26:@14573.4]
  wire  _T_13084; // @[LoadQueue.scala 141:18:@14574.4]
  wire  entriesToCheck_8_13; // @[LoadQueue.scala 141:26:@14575.4]
  wire  _T_13086; // @[LoadQueue.scala 141:18:@14576.4]
  wire  entriesToCheck_8_14; // @[LoadQueue.scala 141:26:@14577.4]
  wire  _T_13088; // @[LoadQueue.scala 141:18:@14578.4]
  wire  entriesToCheck_8_15; // @[LoadQueue.scala 141:26:@14579.4]
  wire  _T_13090; // @[LoadQueue.scala 141:18:@14596.4]
  wire  entriesToCheck_9_0; // @[LoadQueue.scala 141:26:@14597.4]
  wire  _T_13092; // @[LoadQueue.scala 141:18:@14598.4]
  wire  entriesToCheck_9_1; // @[LoadQueue.scala 141:26:@14599.4]
  wire  _T_13094; // @[LoadQueue.scala 141:18:@14600.4]
  wire  entriesToCheck_9_2; // @[LoadQueue.scala 141:26:@14601.4]
  wire  _T_13096; // @[LoadQueue.scala 141:18:@14602.4]
  wire  entriesToCheck_9_3; // @[LoadQueue.scala 141:26:@14603.4]
  wire  _T_13098; // @[LoadQueue.scala 141:18:@14604.4]
  wire  entriesToCheck_9_4; // @[LoadQueue.scala 141:26:@14605.4]
  wire  _T_13100; // @[LoadQueue.scala 141:18:@14606.4]
  wire  entriesToCheck_9_5; // @[LoadQueue.scala 141:26:@14607.4]
  wire  _T_13102; // @[LoadQueue.scala 141:18:@14608.4]
  wire  entriesToCheck_9_6; // @[LoadQueue.scala 141:26:@14609.4]
  wire  _T_13104; // @[LoadQueue.scala 141:18:@14610.4]
  wire  entriesToCheck_9_7; // @[LoadQueue.scala 141:26:@14611.4]
  wire  _T_13106; // @[LoadQueue.scala 141:18:@14612.4]
  wire  entriesToCheck_9_8; // @[LoadQueue.scala 141:26:@14613.4]
  wire  _T_13108; // @[LoadQueue.scala 141:18:@14614.4]
  wire  entriesToCheck_9_9; // @[LoadQueue.scala 141:26:@14615.4]
  wire  _T_13110; // @[LoadQueue.scala 141:18:@14616.4]
  wire  entriesToCheck_9_10; // @[LoadQueue.scala 141:26:@14617.4]
  wire  _T_13112; // @[LoadQueue.scala 141:18:@14618.4]
  wire  entriesToCheck_9_11; // @[LoadQueue.scala 141:26:@14619.4]
  wire  _T_13114; // @[LoadQueue.scala 141:18:@14620.4]
  wire  entriesToCheck_9_12; // @[LoadQueue.scala 141:26:@14621.4]
  wire  _T_13116; // @[LoadQueue.scala 141:18:@14622.4]
  wire  entriesToCheck_9_13; // @[LoadQueue.scala 141:26:@14623.4]
  wire  _T_13118; // @[LoadQueue.scala 141:18:@14624.4]
  wire  entriesToCheck_9_14; // @[LoadQueue.scala 141:26:@14625.4]
  wire  _T_13120; // @[LoadQueue.scala 141:18:@14626.4]
  wire  entriesToCheck_9_15; // @[LoadQueue.scala 141:26:@14627.4]
  wire  _T_13122; // @[LoadQueue.scala 141:18:@14644.4]
  wire  entriesToCheck_10_0; // @[LoadQueue.scala 141:26:@14645.4]
  wire  _T_13124; // @[LoadQueue.scala 141:18:@14646.4]
  wire  entriesToCheck_10_1; // @[LoadQueue.scala 141:26:@14647.4]
  wire  _T_13126; // @[LoadQueue.scala 141:18:@14648.4]
  wire  entriesToCheck_10_2; // @[LoadQueue.scala 141:26:@14649.4]
  wire  _T_13128; // @[LoadQueue.scala 141:18:@14650.4]
  wire  entriesToCheck_10_3; // @[LoadQueue.scala 141:26:@14651.4]
  wire  _T_13130; // @[LoadQueue.scala 141:18:@14652.4]
  wire  entriesToCheck_10_4; // @[LoadQueue.scala 141:26:@14653.4]
  wire  _T_13132; // @[LoadQueue.scala 141:18:@14654.4]
  wire  entriesToCheck_10_5; // @[LoadQueue.scala 141:26:@14655.4]
  wire  _T_13134; // @[LoadQueue.scala 141:18:@14656.4]
  wire  entriesToCheck_10_6; // @[LoadQueue.scala 141:26:@14657.4]
  wire  _T_13136; // @[LoadQueue.scala 141:18:@14658.4]
  wire  entriesToCheck_10_7; // @[LoadQueue.scala 141:26:@14659.4]
  wire  _T_13138; // @[LoadQueue.scala 141:18:@14660.4]
  wire  entriesToCheck_10_8; // @[LoadQueue.scala 141:26:@14661.4]
  wire  _T_13140; // @[LoadQueue.scala 141:18:@14662.4]
  wire  entriesToCheck_10_9; // @[LoadQueue.scala 141:26:@14663.4]
  wire  _T_13142; // @[LoadQueue.scala 141:18:@14664.4]
  wire  entriesToCheck_10_10; // @[LoadQueue.scala 141:26:@14665.4]
  wire  _T_13144; // @[LoadQueue.scala 141:18:@14666.4]
  wire  entriesToCheck_10_11; // @[LoadQueue.scala 141:26:@14667.4]
  wire  _T_13146; // @[LoadQueue.scala 141:18:@14668.4]
  wire  entriesToCheck_10_12; // @[LoadQueue.scala 141:26:@14669.4]
  wire  _T_13148; // @[LoadQueue.scala 141:18:@14670.4]
  wire  entriesToCheck_10_13; // @[LoadQueue.scala 141:26:@14671.4]
  wire  _T_13150; // @[LoadQueue.scala 141:18:@14672.4]
  wire  entriesToCheck_10_14; // @[LoadQueue.scala 141:26:@14673.4]
  wire  _T_13152; // @[LoadQueue.scala 141:18:@14674.4]
  wire  entriesToCheck_10_15; // @[LoadQueue.scala 141:26:@14675.4]
  wire  _T_13154; // @[LoadQueue.scala 141:18:@14692.4]
  wire  entriesToCheck_11_0; // @[LoadQueue.scala 141:26:@14693.4]
  wire  _T_13156; // @[LoadQueue.scala 141:18:@14694.4]
  wire  entriesToCheck_11_1; // @[LoadQueue.scala 141:26:@14695.4]
  wire  _T_13158; // @[LoadQueue.scala 141:18:@14696.4]
  wire  entriesToCheck_11_2; // @[LoadQueue.scala 141:26:@14697.4]
  wire  _T_13160; // @[LoadQueue.scala 141:18:@14698.4]
  wire  entriesToCheck_11_3; // @[LoadQueue.scala 141:26:@14699.4]
  wire  _T_13162; // @[LoadQueue.scala 141:18:@14700.4]
  wire  entriesToCheck_11_4; // @[LoadQueue.scala 141:26:@14701.4]
  wire  _T_13164; // @[LoadQueue.scala 141:18:@14702.4]
  wire  entriesToCheck_11_5; // @[LoadQueue.scala 141:26:@14703.4]
  wire  _T_13166; // @[LoadQueue.scala 141:18:@14704.4]
  wire  entriesToCheck_11_6; // @[LoadQueue.scala 141:26:@14705.4]
  wire  _T_13168; // @[LoadQueue.scala 141:18:@14706.4]
  wire  entriesToCheck_11_7; // @[LoadQueue.scala 141:26:@14707.4]
  wire  _T_13170; // @[LoadQueue.scala 141:18:@14708.4]
  wire  entriesToCheck_11_8; // @[LoadQueue.scala 141:26:@14709.4]
  wire  _T_13172; // @[LoadQueue.scala 141:18:@14710.4]
  wire  entriesToCheck_11_9; // @[LoadQueue.scala 141:26:@14711.4]
  wire  _T_13174; // @[LoadQueue.scala 141:18:@14712.4]
  wire  entriesToCheck_11_10; // @[LoadQueue.scala 141:26:@14713.4]
  wire  _T_13176; // @[LoadQueue.scala 141:18:@14714.4]
  wire  entriesToCheck_11_11; // @[LoadQueue.scala 141:26:@14715.4]
  wire  _T_13178; // @[LoadQueue.scala 141:18:@14716.4]
  wire  entriesToCheck_11_12; // @[LoadQueue.scala 141:26:@14717.4]
  wire  _T_13180; // @[LoadQueue.scala 141:18:@14718.4]
  wire  entriesToCheck_11_13; // @[LoadQueue.scala 141:26:@14719.4]
  wire  _T_13182; // @[LoadQueue.scala 141:18:@14720.4]
  wire  entriesToCheck_11_14; // @[LoadQueue.scala 141:26:@14721.4]
  wire  _T_13184; // @[LoadQueue.scala 141:18:@14722.4]
  wire  entriesToCheck_11_15; // @[LoadQueue.scala 141:26:@14723.4]
  wire  _T_13186; // @[LoadQueue.scala 141:18:@14740.4]
  wire  entriesToCheck_12_0; // @[LoadQueue.scala 141:26:@14741.4]
  wire  _T_13188; // @[LoadQueue.scala 141:18:@14742.4]
  wire  entriesToCheck_12_1; // @[LoadQueue.scala 141:26:@14743.4]
  wire  _T_13190; // @[LoadQueue.scala 141:18:@14744.4]
  wire  entriesToCheck_12_2; // @[LoadQueue.scala 141:26:@14745.4]
  wire  _T_13192; // @[LoadQueue.scala 141:18:@14746.4]
  wire  entriesToCheck_12_3; // @[LoadQueue.scala 141:26:@14747.4]
  wire  _T_13194; // @[LoadQueue.scala 141:18:@14748.4]
  wire  entriesToCheck_12_4; // @[LoadQueue.scala 141:26:@14749.4]
  wire  _T_13196; // @[LoadQueue.scala 141:18:@14750.4]
  wire  entriesToCheck_12_5; // @[LoadQueue.scala 141:26:@14751.4]
  wire  _T_13198; // @[LoadQueue.scala 141:18:@14752.4]
  wire  entriesToCheck_12_6; // @[LoadQueue.scala 141:26:@14753.4]
  wire  _T_13200; // @[LoadQueue.scala 141:18:@14754.4]
  wire  entriesToCheck_12_7; // @[LoadQueue.scala 141:26:@14755.4]
  wire  _T_13202; // @[LoadQueue.scala 141:18:@14756.4]
  wire  entriesToCheck_12_8; // @[LoadQueue.scala 141:26:@14757.4]
  wire  _T_13204; // @[LoadQueue.scala 141:18:@14758.4]
  wire  entriesToCheck_12_9; // @[LoadQueue.scala 141:26:@14759.4]
  wire  _T_13206; // @[LoadQueue.scala 141:18:@14760.4]
  wire  entriesToCheck_12_10; // @[LoadQueue.scala 141:26:@14761.4]
  wire  _T_13208; // @[LoadQueue.scala 141:18:@14762.4]
  wire  entriesToCheck_12_11; // @[LoadQueue.scala 141:26:@14763.4]
  wire  _T_13210; // @[LoadQueue.scala 141:18:@14764.4]
  wire  entriesToCheck_12_12; // @[LoadQueue.scala 141:26:@14765.4]
  wire  _T_13212; // @[LoadQueue.scala 141:18:@14766.4]
  wire  entriesToCheck_12_13; // @[LoadQueue.scala 141:26:@14767.4]
  wire  _T_13214; // @[LoadQueue.scala 141:18:@14768.4]
  wire  entriesToCheck_12_14; // @[LoadQueue.scala 141:26:@14769.4]
  wire  _T_13216; // @[LoadQueue.scala 141:18:@14770.4]
  wire  entriesToCheck_12_15; // @[LoadQueue.scala 141:26:@14771.4]
  wire  _T_13218; // @[LoadQueue.scala 141:18:@14788.4]
  wire  entriesToCheck_13_0; // @[LoadQueue.scala 141:26:@14789.4]
  wire  _T_13220; // @[LoadQueue.scala 141:18:@14790.4]
  wire  entriesToCheck_13_1; // @[LoadQueue.scala 141:26:@14791.4]
  wire  _T_13222; // @[LoadQueue.scala 141:18:@14792.4]
  wire  entriesToCheck_13_2; // @[LoadQueue.scala 141:26:@14793.4]
  wire  _T_13224; // @[LoadQueue.scala 141:18:@14794.4]
  wire  entriesToCheck_13_3; // @[LoadQueue.scala 141:26:@14795.4]
  wire  _T_13226; // @[LoadQueue.scala 141:18:@14796.4]
  wire  entriesToCheck_13_4; // @[LoadQueue.scala 141:26:@14797.4]
  wire  _T_13228; // @[LoadQueue.scala 141:18:@14798.4]
  wire  entriesToCheck_13_5; // @[LoadQueue.scala 141:26:@14799.4]
  wire  _T_13230; // @[LoadQueue.scala 141:18:@14800.4]
  wire  entriesToCheck_13_6; // @[LoadQueue.scala 141:26:@14801.4]
  wire  _T_13232; // @[LoadQueue.scala 141:18:@14802.4]
  wire  entriesToCheck_13_7; // @[LoadQueue.scala 141:26:@14803.4]
  wire  _T_13234; // @[LoadQueue.scala 141:18:@14804.4]
  wire  entriesToCheck_13_8; // @[LoadQueue.scala 141:26:@14805.4]
  wire  _T_13236; // @[LoadQueue.scala 141:18:@14806.4]
  wire  entriesToCheck_13_9; // @[LoadQueue.scala 141:26:@14807.4]
  wire  _T_13238; // @[LoadQueue.scala 141:18:@14808.4]
  wire  entriesToCheck_13_10; // @[LoadQueue.scala 141:26:@14809.4]
  wire  _T_13240; // @[LoadQueue.scala 141:18:@14810.4]
  wire  entriesToCheck_13_11; // @[LoadQueue.scala 141:26:@14811.4]
  wire  _T_13242; // @[LoadQueue.scala 141:18:@14812.4]
  wire  entriesToCheck_13_12; // @[LoadQueue.scala 141:26:@14813.4]
  wire  _T_13244; // @[LoadQueue.scala 141:18:@14814.4]
  wire  entriesToCheck_13_13; // @[LoadQueue.scala 141:26:@14815.4]
  wire  _T_13246; // @[LoadQueue.scala 141:18:@14816.4]
  wire  entriesToCheck_13_14; // @[LoadQueue.scala 141:26:@14817.4]
  wire  _T_13248; // @[LoadQueue.scala 141:18:@14818.4]
  wire  entriesToCheck_13_15; // @[LoadQueue.scala 141:26:@14819.4]
  wire  _T_13250; // @[LoadQueue.scala 141:18:@14836.4]
  wire  entriesToCheck_14_0; // @[LoadQueue.scala 141:26:@14837.4]
  wire  _T_13252; // @[LoadQueue.scala 141:18:@14838.4]
  wire  entriesToCheck_14_1; // @[LoadQueue.scala 141:26:@14839.4]
  wire  _T_13254; // @[LoadQueue.scala 141:18:@14840.4]
  wire  entriesToCheck_14_2; // @[LoadQueue.scala 141:26:@14841.4]
  wire  _T_13256; // @[LoadQueue.scala 141:18:@14842.4]
  wire  entriesToCheck_14_3; // @[LoadQueue.scala 141:26:@14843.4]
  wire  _T_13258; // @[LoadQueue.scala 141:18:@14844.4]
  wire  entriesToCheck_14_4; // @[LoadQueue.scala 141:26:@14845.4]
  wire  _T_13260; // @[LoadQueue.scala 141:18:@14846.4]
  wire  entriesToCheck_14_5; // @[LoadQueue.scala 141:26:@14847.4]
  wire  _T_13262; // @[LoadQueue.scala 141:18:@14848.4]
  wire  entriesToCheck_14_6; // @[LoadQueue.scala 141:26:@14849.4]
  wire  _T_13264; // @[LoadQueue.scala 141:18:@14850.4]
  wire  entriesToCheck_14_7; // @[LoadQueue.scala 141:26:@14851.4]
  wire  _T_13266; // @[LoadQueue.scala 141:18:@14852.4]
  wire  entriesToCheck_14_8; // @[LoadQueue.scala 141:26:@14853.4]
  wire  _T_13268; // @[LoadQueue.scala 141:18:@14854.4]
  wire  entriesToCheck_14_9; // @[LoadQueue.scala 141:26:@14855.4]
  wire  _T_13270; // @[LoadQueue.scala 141:18:@14856.4]
  wire  entriesToCheck_14_10; // @[LoadQueue.scala 141:26:@14857.4]
  wire  _T_13272; // @[LoadQueue.scala 141:18:@14858.4]
  wire  entriesToCheck_14_11; // @[LoadQueue.scala 141:26:@14859.4]
  wire  _T_13274; // @[LoadQueue.scala 141:18:@14860.4]
  wire  entriesToCheck_14_12; // @[LoadQueue.scala 141:26:@14861.4]
  wire  _T_13276; // @[LoadQueue.scala 141:18:@14862.4]
  wire  entriesToCheck_14_13; // @[LoadQueue.scala 141:26:@14863.4]
  wire  _T_13278; // @[LoadQueue.scala 141:18:@14864.4]
  wire  entriesToCheck_14_14; // @[LoadQueue.scala 141:26:@14865.4]
  wire  _T_13280; // @[LoadQueue.scala 141:18:@14866.4]
  wire  entriesToCheck_14_15; // @[LoadQueue.scala 141:26:@14867.4]
  wire  _T_13282; // @[LoadQueue.scala 141:18:@14884.4]
  wire  entriesToCheck_15_0; // @[LoadQueue.scala 141:26:@14885.4]
  wire  _T_13284; // @[LoadQueue.scala 141:18:@14886.4]
  wire  entriesToCheck_15_1; // @[LoadQueue.scala 141:26:@14887.4]
  wire  _T_13286; // @[LoadQueue.scala 141:18:@14888.4]
  wire  entriesToCheck_15_2; // @[LoadQueue.scala 141:26:@14889.4]
  wire  _T_13288; // @[LoadQueue.scala 141:18:@14890.4]
  wire  entriesToCheck_15_3; // @[LoadQueue.scala 141:26:@14891.4]
  wire  _T_13290; // @[LoadQueue.scala 141:18:@14892.4]
  wire  entriesToCheck_15_4; // @[LoadQueue.scala 141:26:@14893.4]
  wire  _T_13292; // @[LoadQueue.scala 141:18:@14894.4]
  wire  entriesToCheck_15_5; // @[LoadQueue.scala 141:26:@14895.4]
  wire  _T_13294; // @[LoadQueue.scala 141:18:@14896.4]
  wire  entriesToCheck_15_6; // @[LoadQueue.scala 141:26:@14897.4]
  wire  _T_13296; // @[LoadQueue.scala 141:18:@14898.4]
  wire  entriesToCheck_15_7; // @[LoadQueue.scala 141:26:@14899.4]
  wire  _T_13298; // @[LoadQueue.scala 141:18:@14900.4]
  wire  entriesToCheck_15_8; // @[LoadQueue.scala 141:26:@14901.4]
  wire  _T_13300; // @[LoadQueue.scala 141:18:@14902.4]
  wire  entriesToCheck_15_9; // @[LoadQueue.scala 141:26:@14903.4]
  wire  _T_13302; // @[LoadQueue.scala 141:18:@14904.4]
  wire  entriesToCheck_15_10; // @[LoadQueue.scala 141:26:@14905.4]
  wire  _T_13304; // @[LoadQueue.scala 141:18:@14906.4]
  wire  entriesToCheck_15_11; // @[LoadQueue.scala 141:26:@14907.4]
  wire  _T_13306; // @[LoadQueue.scala 141:18:@14908.4]
  wire  entriesToCheck_15_12; // @[LoadQueue.scala 141:26:@14909.4]
  wire  _T_13308; // @[LoadQueue.scala 141:18:@14910.4]
  wire  entriesToCheck_15_13; // @[LoadQueue.scala 141:26:@14911.4]
  wire  _T_13310; // @[LoadQueue.scala 141:18:@14912.4]
  wire  entriesToCheck_15_14; // @[LoadQueue.scala 141:26:@14913.4]
  wire  _T_13312; // @[LoadQueue.scala 141:18:@14914.4]
  wire  entriesToCheck_15_15; // @[LoadQueue.scala 141:26:@14915.4]
  wire  _T_14544; // @[LoadQueue.scala 151:92:@14933.4]
  wire  _T_14545; // @[LoadQueue.scala 152:41:@14934.4]
  wire  _T_14546; // @[LoadQueue.scala 153:30:@14935.4]
  wire  conflict_0_0; // @[LoadQueue.scala 152:68:@14936.4]
  wire  _T_14548; // @[LoadQueue.scala 151:92:@14938.4]
  wire  _T_14549; // @[LoadQueue.scala 152:41:@14939.4]
  wire  _T_14550; // @[LoadQueue.scala 153:30:@14940.4]
  wire  conflict_0_1; // @[LoadQueue.scala 152:68:@14941.4]
  wire  _T_14552; // @[LoadQueue.scala 151:92:@14943.4]
  wire  _T_14553; // @[LoadQueue.scala 152:41:@14944.4]
  wire  _T_14554; // @[LoadQueue.scala 153:30:@14945.4]
  wire  conflict_0_2; // @[LoadQueue.scala 152:68:@14946.4]
  wire  _T_14556; // @[LoadQueue.scala 151:92:@14948.4]
  wire  _T_14557; // @[LoadQueue.scala 152:41:@14949.4]
  wire  _T_14558; // @[LoadQueue.scala 153:30:@14950.4]
  wire  conflict_0_3; // @[LoadQueue.scala 152:68:@14951.4]
  wire  _T_14560; // @[LoadQueue.scala 151:92:@14953.4]
  wire  _T_14561; // @[LoadQueue.scala 152:41:@14954.4]
  wire  _T_14562; // @[LoadQueue.scala 153:30:@14955.4]
  wire  conflict_0_4; // @[LoadQueue.scala 152:68:@14956.4]
  wire  _T_14564; // @[LoadQueue.scala 151:92:@14958.4]
  wire  _T_14565; // @[LoadQueue.scala 152:41:@14959.4]
  wire  _T_14566; // @[LoadQueue.scala 153:30:@14960.4]
  wire  conflict_0_5; // @[LoadQueue.scala 152:68:@14961.4]
  wire  _T_14568; // @[LoadQueue.scala 151:92:@14963.4]
  wire  _T_14569; // @[LoadQueue.scala 152:41:@14964.4]
  wire  _T_14570; // @[LoadQueue.scala 153:30:@14965.4]
  wire  conflict_0_6; // @[LoadQueue.scala 152:68:@14966.4]
  wire  _T_14572; // @[LoadQueue.scala 151:92:@14968.4]
  wire  _T_14573; // @[LoadQueue.scala 152:41:@14969.4]
  wire  _T_14574; // @[LoadQueue.scala 153:30:@14970.4]
  wire  conflict_0_7; // @[LoadQueue.scala 152:68:@14971.4]
  wire  _T_14576; // @[LoadQueue.scala 151:92:@14973.4]
  wire  _T_14577; // @[LoadQueue.scala 152:41:@14974.4]
  wire  _T_14578; // @[LoadQueue.scala 153:30:@14975.4]
  wire  conflict_0_8; // @[LoadQueue.scala 152:68:@14976.4]
  wire  _T_14580; // @[LoadQueue.scala 151:92:@14978.4]
  wire  _T_14581; // @[LoadQueue.scala 152:41:@14979.4]
  wire  _T_14582; // @[LoadQueue.scala 153:30:@14980.4]
  wire  conflict_0_9; // @[LoadQueue.scala 152:68:@14981.4]
  wire  _T_14584; // @[LoadQueue.scala 151:92:@14983.4]
  wire  _T_14585; // @[LoadQueue.scala 152:41:@14984.4]
  wire  _T_14586; // @[LoadQueue.scala 153:30:@14985.4]
  wire  conflict_0_10; // @[LoadQueue.scala 152:68:@14986.4]
  wire  _T_14588; // @[LoadQueue.scala 151:92:@14988.4]
  wire  _T_14589; // @[LoadQueue.scala 152:41:@14989.4]
  wire  _T_14590; // @[LoadQueue.scala 153:30:@14990.4]
  wire  conflict_0_11; // @[LoadQueue.scala 152:68:@14991.4]
  wire  _T_14592; // @[LoadQueue.scala 151:92:@14993.4]
  wire  _T_14593; // @[LoadQueue.scala 152:41:@14994.4]
  wire  _T_14594; // @[LoadQueue.scala 153:30:@14995.4]
  wire  conflict_0_12; // @[LoadQueue.scala 152:68:@14996.4]
  wire  _T_14596; // @[LoadQueue.scala 151:92:@14998.4]
  wire  _T_14597; // @[LoadQueue.scala 152:41:@14999.4]
  wire  _T_14598; // @[LoadQueue.scala 153:30:@15000.4]
  wire  conflict_0_13; // @[LoadQueue.scala 152:68:@15001.4]
  wire  _T_14600; // @[LoadQueue.scala 151:92:@15003.4]
  wire  _T_14601; // @[LoadQueue.scala 152:41:@15004.4]
  wire  _T_14602; // @[LoadQueue.scala 153:30:@15005.4]
  wire  conflict_0_14; // @[LoadQueue.scala 152:68:@15006.4]
  wire  _T_14604; // @[LoadQueue.scala 151:92:@15008.4]
  wire  _T_14605; // @[LoadQueue.scala 152:41:@15009.4]
  wire  _T_14606; // @[LoadQueue.scala 153:30:@15010.4]
  wire  conflict_0_15; // @[LoadQueue.scala 152:68:@15011.4]
  wire  _T_14608; // @[LoadQueue.scala 151:92:@15013.4]
  wire  _T_14609; // @[LoadQueue.scala 152:41:@15014.4]
  wire  _T_14610; // @[LoadQueue.scala 153:30:@15015.4]
  wire  conflict_1_0; // @[LoadQueue.scala 152:68:@15016.4]
  wire  _T_14612; // @[LoadQueue.scala 151:92:@15018.4]
  wire  _T_14613; // @[LoadQueue.scala 152:41:@15019.4]
  wire  _T_14614; // @[LoadQueue.scala 153:30:@15020.4]
  wire  conflict_1_1; // @[LoadQueue.scala 152:68:@15021.4]
  wire  _T_14616; // @[LoadQueue.scala 151:92:@15023.4]
  wire  _T_14617; // @[LoadQueue.scala 152:41:@15024.4]
  wire  _T_14618; // @[LoadQueue.scala 153:30:@15025.4]
  wire  conflict_1_2; // @[LoadQueue.scala 152:68:@15026.4]
  wire  _T_14620; // @[LoadQueue.scala 151:92:@15028.4]
  wire  _T_14621; // @[LoadQueue.scala 152:41:@15029.4]
  wire  _T_14622; // @[LoadQueue.scala 153:30:@15030.4]
  wire  conflict_1_3; // @[LoadQueue.scala 152:68:@15031.4]
  wire  _T_14624; // @[LoadQueue.scala 151:92:@15033.4]
  wire  _T_14625; // @[LoadQueue.scala 152:41:@15034.4]
  wire  _T_14626; // @[LoadQueue.scala 153:30:@15035.4]
  wire  conflict_1_4; // @[LoadQueue.scala 152:68:@15036.4]
  wire  _T_14628; // @[LoadQueue.scala 151:92:@15038.4]
  wire  _T_14629; // @[LoadQueue.scala 152:41:@15039.4]
  wire  _T_14630; // @[LoadQueue.scala 153:30:@15040.4]
  wire  conflict_1_5; // @[LoadQueue.scala 152:68:@15041.4]
  wire  _T_14632; // @[LoadQueue.scala 151:92:@15043.4]
  wire  _T_14633; // @[LoadQueue.scala 152:41:@15044.4]
  wire  _T_14634; // @[LoadQueue.scala 153:30:@15045.4]
  wire  conflict_1_6; // @[LoadQueue.scala 152:68:@15046.4]
  wire  _T_14636; // @[LoadQueue.scala 151:92:@15048.4]
  wire  _T_14637; // @[LoadQueue.scala 152:41:@15049.4]
  wire  _T_14638; // @[LoadQueue.scala 153:30:@15050.4]
  wire  conflict_1_7; // @[LoadQueue.scala 152:68:@15051.4]
  wire  _T_14640; // @[LoadQueue.scala 151:92:@15053.4]
  wire  _T_14641; // @[LoadQueue.scala 152:41:@15054.4]
  wire  _T_14642; // @[LoadQueue.scala 153:30:@15055.4]
  wire  conflict_1_8; // @[LoadQueue.scala 152:68:@15056.4]
  wire  _T_14644; // @[LoadQueue.scala 151:92:@15058.4]
  wire  _T_14645; // @[LoadQueue.scala 152:41:@15059.4]
  wire  _T_14646; // @[LoadQueue.scala 153:30:@15060.4]
  wire  conflict_1_9; // @[LoadQueue.scala 152:68:@15061.4]
  wire  _T_14648; // @[LoadQueue.scala 151:92:@15063.4]
  wire  _T_14649; // @[LoadQueue.scala 152:41:@15064.4]
  wire  _T_14650; // @[LoadQueue.scala 153:30:@15065.4]
  wire  conflict_1_10; // @[LoadQueue.scala 152:68:@15066.4]
  wire  _T_14652; // @[LoadQueue.scala 151:92:@15068.4]
  wire  _T_14653; // @[LoadQueue.scala 152:41:@15069.4]
  wire  _T_14654; // @[LoadQueue.scala 153:30:@15070.4]
  wire  conflict_1_11; // @[LoadQueue.scala 152:68:@15071.4]
  wire  _T_14656; // @[LoadQueue.scala 151:92:@15073.4]
  wire  _T_14657; // @[LoadQueue.scala 152:41:@15074.4]
  wire  _T_14658; // @[LoadQueue.scala 153:30:@15075.4]
  wire  conflict_1_12; // @[LoadQueue.scala 152:68:@15076.4]
  wire  _T_14660; // @[LoadQueue.scala 151:92:@15078.4]
  wire  _T_14661; // @[LoadQueue.scala 152:41:@15079.4]
  wire  _T_14662; // @[LoadQueue.scala 153:30:@15080.4]
  wire  conflict_1_13; // @[LoadQueue.scala 152:68:@15081.4]
  wire  _T_14664; // @[LoadQueue.scala 151:92:@15083.4]
  wire  _T_14665; // @[LoadQueue.scala 152:41:@15084.4]
  wire  _T_14666; // @[LoadQueue.scala 153:30:@15085.4]
  wire  conflict_1_14; // @[LoadQueue.scala 152:68:@15086.4]
  wire  _T_14668; // @[LoadQueue.scala 151:92:@15088.4]
  wire  _T_14669; // @[LoadQueue.scala 152:41:@15089.4]
  wire  _T_14670; // @[LoadQueue.scala 153:30:@15090.4]
  wire  conflict_1_15; // @[LoadQueue.scala 152:68:@15091.4]
  wire  _T_14672; // @[LoadQueue.scala 151:92:@15093.4]
  wire  _T_14673; // @[LoadQueue.scala 152:41:@15094.4]
  wire  _T_14674; // @[LoadQueue.scala 153:30:@15095.4]
  wire  conflict_2_0; // @[LoadQueue.scala 152:68:@15096.4]
  wire  _T_14676; // @[LoadQueue.scala 151:92:@15098.4]
  wire  _T_14677; // @[LoadQueue.scala 152:41:@15099.4]
  wire  _T_14678; // @[LoadQueue.scala 153:30:@15100.4]
  wire  conflict_2_1; // @[LoadQueue.scala 152:68:@15101.4]
  wire  _T_14680; // @[LoadQueue.scala 151:92:@15103.4]
  wire  _T_14681; // @[LoadQueue.scala 152:41:@15104.4]
  wire  _T_14682; // @[LoadQueue.scala 153:30:@15105.4]
  wire  conflict_2_2; // @[LoadQueue.scala 152:68:@15106.4]
  wire  _T_14684; // @[LoadQueue.scala 151:92:@15108.4]
  wire  _T_14685; // @[LoadQueue.scala 152:41:@15109.4]
  wire  _T_14686; // @[LoadQueue.scala 153:30:@15110.4]
  wire  conflict_2_3; // @[LoadQueue.scala 152:68:@15111.4]
  wire  _T_14688; // @[LoadQueue.scala 151:92:@15113.4]
  wire  _T_14689; // @[LoadQueue.scala 152:41:@15114.4]
  wire  _T_14690; // @[LoadQueue.scala 153:30:@15115.4]
  wire  conflict_2_4; // @[LoadQueue.scala 152:68:@15116.4]
  wire  _T_14692; // @[LoadQueue.scala 151:92:@15118.4]
  wire  _T_14693; // @[LoadQueue.scala 152:41:@15119.4]
  wire  _T_14694; // @[LoadQueue.scala 153:30:@15120.4]
  wire  conflict_2_5; // @[LoadQueue.scala 152:68:@15121.4]
  wire  _T_14696; // @[LoadQueue.scala 151:92:@15123.4]
  wire  _T_14697; // @[LoadQueue.scala 152:41:@15124.4]
  wire  _T_14698; // @[LoadQueue.scala 153:30:@15125.4]
  wire  conflict_2_6; // @[LoadQueue.scala 152:68:@15126.4]
  wire  _T_14700; // @[LoadQueue.scala 151:92:@15128.4]
  wire  _T_14701; // @[LoadQueue.scala 152:41:@15129.4]
  wire  _T_14702; // @[LoadQueue.scala 153:30:@15130.4]
  wire  conflict_2_7; // @[LoadQueue.scala 152:68:@15131.4]
  wire  _T_14704; // @[LoadQueue.scala 151:92:@15133.4]
  wire  _T_14705; // @[LoadQueue.scala 152:41:@15134.4]
  wire  _T_14706; // @[LoadQueue.scala 153:30:@15135.4]
  wire  conflict_2_8; // @[LoadQueue.scala 152:68:@15136.4]
  wire  _T_14708; // @[LoadQueue.scala 151:92:@15138.4]
  wire  _T_14709; // @[LoadQueue.scala 152:41:@15139.4]
  wire  _T_14710; // @[LoadQueue.scala 153:30:@15140.4]
  wire  conflict_2_9; // @[LoadQueue.scala 152:68:@15141.4]
  wire  _T_14712; // @[LoadQueue.scala 151:92:@15143.4]
  wire  _T_14713; // @[LoadQueue.scala 152:41:@15144.4]
  wire  _T_14714; // @[LoadQueue.scala 153:30:@15145.4]
  wire  conflict_2_10; // @[LoadQueue.scala 152:68:@15146.4]
  wire  _T_14716; // @[LoadQueue.scala 151:92:@15148.4]
  wire  _T_14717; // @[LoadQueue.scala 152:41:@15149.4]
  wire  _T_14718; // @[LoadQueue.scala 153:30:@15150.4]
  wire  conflict_2_11; // @[LoadQueue.scala 152:68:@15151.4]
  wire  _T_14720; // @[LoadQueue.scala 151:92:@15153.4]
  wire  _T_14721; // @[LoadQueue.scala 152:41:@15154.4]
  wire  _T_14722; // @[LoadQueue.scala 153:30:@15155.4]
  wire  conflict_2_12; // @[LoadQueue.scala 152:68:@15156.4]
  wire  _T_14724; // @[LoadQueue.scala 151:92:@15158.4]
  wire  _T_14725; // @[LoadQueue.scala 152:41:@15159.4]
  wire  _T_14726; // @[LoadQueue.scala 153:30:@15160.4]
  wire  conflict_2_13; // @[LoadQueue.scala 152:68:@15161.4]
  wire  _T_14728; // @[LoadQueue.scala 151:92:@15163.4]
  wire  _T_14729; // @[LoadQueue.scala 152:41:@15164.4]
  wire  _T_14730; // @[LoadQueue.scala 153:30:@15165.4]
  wire  conflict_2_14; // @[LoadQueue.scala 152:68:@15166.4]
  wire  _T_14732; // @[LoadQueue.scala 151:92:@15168.4]
  wire  _T_14733; // @[LoadQueue.scala 152:41:@15169.4]
  wire  _T_14734; // @[LoadQueue.scala 153:30:@15170.4]
  wire  conflict_2_15; // @[LoadQueue.scala 152:68:@15171.4]
  wire  _T_14736; // @[LoadQueue.scala 151:92:@15173.4]
  wire  _T_14737; // @[LoadQueue.scala 152:41:@15174.4]
  wire  _T_14738; // @[LoadQueue.scala 153:30:@15175.4]
  wire  conflict_3_0; // @[LoadQueue.scala 152:68:@15176.4]
  wire  _T_14740; // @[LoadQueue.scala 151:92:@15178.4]
  wire  _T_14741; // @[LoadQueue.scala 152:41:@15179.4]
  wire  _T_14742; // @[LoadQueue.scala 153:30:@15180.4]
  wire  conflict_3_1; // @[LoadQueue.scala 152:68:@15181.4]
  wire  _T_14744; // @[LoadQueue.scala 151:92:@15183.4]
  wire  _T_14745; // @[LoadQueue.scala 152:41:@15184.4]
  wire  _T_14746; // @[LoadQueue.scala 153:30:@15185.4]
  wire  conflict_3_2; // @[LoadQueue.scala 152:68:@15186.4]
  wire  _T_14748; // @[LoadQueue.scala 151:92:@15188.4]
  wire  _T_14749; // @[LoadQueue.scala 152:41:@15189.4]
  wire  _T_14750; // @[LoadQueue.scala 153:30:@15190.4]
  wire  conflict_3_3; // @[LoadQueue.scala 152:68:@15191.4]
  wire  _T_14752; // @[LoadQueue.scala 151:92:@15193.4]
  wire  _T_14753; // @[LoadQueue.scala 152:41:@15194.4]
  wire  _T_14754; // @[LoadQueue.scala 153:30:@15195.4]
  wire  conflict_3_4; // @[LoadQueue.scala 152:68:@15196.4]
  wire  _T_14756; // @[LoadQueue.scala 151:92:@15198.4]
  wire  _T_14757; // @[LoadQueue.scala 152:41:@15199.4]
  wire  _T_14758; // @[LoadQueue.scala 153:30:@15200.4]
  wire  conflict_3_5; // @[LoadQueue.scala 152:68:@15201.4]
  wire  _T_14760; // @[LoadQueue.scala 151:92:@15203.4]
  wire  _T_14761; // @[LoadQueue.scala 152:41:@15204.4]
  wire  _T_14762; // @[LoadQueue.scala 153:30:@15205.4]
  wire  conflict_3_6; // @[LoadQueue.scala 152:68:@15206.4]
  wire  _T_14764; // @[LoadQueue.scala 151:92:@15208.4]
  wire  _T_14765; // @[LoadQueue.scala 152:41:@15209.4]
  wire  _T_14766; // @[LoadQueue.scala 153:30:@15210.4]
  wire  conflict_3_7; // @[LoadQueue.scala 152:68:@15211.4]
  wire  _T_14768; // @[LoadQueue.scala 151:92:@15213.4]
  wire  _T_14769; // @[LoadQueue.scala 152:41:@15214.4]
  wire  _T_14770; // @[LoadQueue.scala 153:30:@15215.4]
  wire  conflict_3_8; // @[LoadQueue.scala 152:68:@15216.4]
  wire  _T_14772; // @[LoadQueue.scala 151:92:@15218.4]
  wire  _T_14773; // @[LoadQueue.scala 152:41:@15219.4]
  wire  _T_14774; // @[LoadQueue.scala 153:30:@15220.4]
  wire  conflict_3_9; // @[LoadQueue.scala 152:68:@15221.4]
  wire  _T_14776; // @[LoadQueue.scala 151:92:@15223.4]
  wire  _T_14777; // @[LoadQueue.scala 152:41:@15224.4]
  wire  _T_14778; // @[LoadQueue.scala 153:30:@15225.4]
  wire  conflict_3_10; // @[LoadQueue.scala 152:68:@15226.4]
  wire  _T_14780; // @[LoadQueue.scala 151:92:@15228.4]
  wire  _T_14781; // @[LoadQueue.scala 152:41:@15229.4]
  wire  _T_14782; // @[LoadQueue.scala 153:30:@15230.4]
  wire  conflict_3_11; // @[LoadQueue.scala 152:68:@15231.4]
  wire  _T_14784; // @[LoadQueue.scala 151:92:@15233.4]
  wire  _T_14785; // @[LoadQueue.scala 152:41:@15234.4]
  wire  _T_14786; // @[LoadQueue.scala 153:30:@15235.4]
  wire  conflict_3_12; // @[LoadQueue.scala 152:68:@15236.4]
  wire  _T_14788; // @[LoadQueue.scala 151:92:@15238.4]
  wire  _T_14789; // @[LoadQueue.scala 152:41:@15239.4]
  wire  _T_14790; // @[LoadQueue.scala 153:30:@15240.4]
  wire  conflict_3_13; // @[LoadQueue.scala 152:68:@15241.4]
  wire  _T_14792; // @[LoadQueue.scala 151:92:@15243.4]
  wire  _T_14793; // @[LoadQueue.scala 152:41:@15244.4]
  wire  _T_14794; // @[LoadQueue.scala 153:30:@15245.4]
  wire  conflict_3_14; // @[LoadQueue.scala 152:68:@15246.4]
  wire  _T_14796; // @[LoadQueue.scala 151:92:@15248.4]
  wire  _T_14797; // @[LoadQueue.scala 152:41:@15249.4]
  wire  _T_14798; // @[LoadQueue.scala 153:30:@15250.4]
  wire  conflict_3_15; // @[LoadQueue.scala 152:68:@15251.4]
  wire  _T_14800; // @[LoadQueue.scala 151:92:@15253.4]
  wire  _T_14801; // @[LoadQueue.scala 152:41:@15254.4]
  wire  _T_14802; // @[LoadQueue.scala 153:30:@15255.4]
  wire  conflict_4_0; // @[LoadQueue.scala 152:68:@15256.4]
  wire  _T_14804; // @[LoadQueue.scala 151:92:@15258.4]
  wire  _T_14805; // @[LoadQueue.scala 152:41:@15259.4]
  wire  _T_14806; // @[LoadQueue.scala 153:30:@15260.4]
  wire  conflict_4_1; // @[LoadQueue.scala 152:68:@15261.4]
  wire  _T_14808; // @[LoadQueue.scala 151:92:@15263.4]
  wire  _T_14809; // @[LoadQueue.scala 152:41:@15264.4]
  wire  _T_14810; // @[LoadQueue.scala 153:30:@15265.4]
  wire  conflict_4_2; // @[LoadQueue.scala 152:68:@15266.4]
  wire  _T_14812; // @[LoadQueue.scala 151:92:@15268.4]
  wire  _T_14813; // @[LoadQueue.scala 152:41:@15269.4]
  wire  _T_14814; // @[LoadQueue.scala 153:30:@15270.4]
  wire  conflict_4_3; // @[LoadQueue.scala 152:68:@15271.4]
  wire  _T_14816; // @[LoadQueue.scala 151:92:@15273.4]
  wire  _T_14817; // @[LoadQueue.scala 152:41:@15274.4]
  wire  _T_14818; // @[LoadQueue.scala 153:30:@15275.4]
  wire  conflict_4_4; // @[LoadQueue.scala 152:68:@15276.4]
  wire  _T_14820; // @[LoadQueue.scala 151:92:@15278.4]
  wire  _T_14821; // @[LoadQueue.scala 152:41:@15279.4]
  wire  _T_14822; // @[LoadQueue.scala 153:30:@15280.4]
  wire  conflict_4_5; // @[LoadQueue.scala 152:68:@15281.4]
  wire  _T_14824; // @[LoadQueue.scala 151:92:@15283.4]
  wire  _T_14825; // @[LoadQueue.scala 152:41:@15284.4]
  wire  _T_14826; // @[LoadQueue.scala 153:30:@15285.4]
  wire  conflict_4_6; // @[LoadQueue.scala 152:68:@15286.4]
  wire  _T_14828; // @[LoadQueue.scala 151:92:@15288.4]
  wire  _T_14829; // @[LoadQueue.scala 152:41:@15289.4]
  wire  _T_14830; // @[LoadQueue.scala 153:30:@15290.4]
  wire  conflict_4_7; // @[LoadQueue.scala 152:68:@15291.4]
  wire  _T_14832; // @[LoadQueue.scala 151:92:@15293.4]
  wire  _T_14833; // @[LoadQueue.scala 152:41:@15294.4]
  wire  _T_14834; // @[LoadQueue.scala 153:30:@15295.4]
  wire  conflict_4_8; // @[LoadQueue.scala 152:68:@15296.4]
  wire  _T_14836; // @[LoadQueue.scala 151:92:@15298.4]
  wire  _T_14837; // @[LoadQueue.scala 152:41:@15299.4]
  wire  _T_14838; // @[LoadQueue.scala 153:30:@15300.4]
  wire  conflict_4_9; // @[LoadQueue.scala 152:68:@15301.4]
  wire  _T_14840; // @[LoadQueue.scala 151:92:@15303.4]
  wire  _T_14841; // @[LoadQueue.scala 152:41:@15304.4]
  wire  _T_14842; // @[LoadQueue.scala 153:30:@15305.4]
  wire  conflict_4_10; // @[LoadQueue.scala 152:68:@15306.4]
  wire  _T_14844; // @[LoadQueue.scala 151:92:@15308.4]
  wire  _T_14845; // @[LoadQueue.scala 152:41:@15309.4]
  wire  _T_14846; // @[LoadQueue.scala 153:30:@15310.4]
  wire  conflict_4_11; // @[LoadQueue.scala 152:68:@15311.4]
  wire  _T_14848; // @[LoadQueue.scala 151:92:@15313.4]
  wire  _T_14849; // @[LoadQueue.scala 152:41:@15314.4]
  wire  _T_14850; // @[LoadQueue.scala 153:30:@15315.4]
  wire  conflict_4_12; // @[LoadQueue.scala 152:68:@15316.4]
  wire  _T_14852; // @[LoadQueue.scala 151:92:@15318.4]
  wire  _T_14853; // @[LoadQueue.scala 152:41:@15319.4]
  wire  _T_14854; // @[LoadQueue.scala 153:30:@15320.4]
  wire  conflict_4_13; // @[LoadQueue.scala 152:68:@15321.4]
  wire  _T_14856; // @[LoadQueue.scala 151:92:@15323.4]
  wire  _T_14857; // @[LoadQueue.scala 152:41:@15324.4]
  wire  _T_14858; // @[LoadQueue.scala 153:30:@15325.4]
  wire  conflict_4_14; // @[LoadQueue.scala 152:68:@15326.4]
  wire  _T_14860; // @[LoadQueue.scala 151:92:@15328.4]
  wire  _T_14861; // @[LoadQueue.scala 152:41:@15329.4]
  wire  _T_14862; // @[LoadQueue.scala 153:30:@15330.4]
  wire  conflict_4_15; // @[LoadQueue.scala 152:68:@15331.4]
  wire  _T_14864; // @[LoadQueue.scala 151:92:@15333.4]
  wire  _T_14865; // @[LoadQueue.scala 152:41:@15334.4]
  wire  _T_14866; // @[LoadQueue.scala 153:30:@15335.4]
  wire  conflict_5_0; // @[LoadQueue.scala 152:68:@15336.4]
  wire  _T_14868; // @[LoadQueue.scala 151:92:@15338.4]
  wire  _T_14869; // @[LoadQueue.scala 152:41:@15339.4]
  wire  _T_14870; // @[LoadQueue.scala 153:30:@15340.4]
  wire  conflict_5_1; // @[LoadQueue.scala 152:68:@15341.4]
  wire  _T_14872; // @[LoadQueue.scala 151:92:@15343.4]
  wire  _T_14873; // @[LoadQueue.scala 152:41:@15344.4]
  wire  _T_14874; // @[LoadQueue.scala 153:30:@15345.4]
  wire  conflict_5_2; // @[LoadQueue.scala 152:68:@15346.4]
  wire  _T_14876; // @[LoadQueue.scala 151:92:@15348.4]
  wire  _T_14877; // @[LoadQueue.scala 152:41:@15349.4]
  wire  _T_14878; // @[LoadQueue.scala 153:30:@15350.4]
  wire  conflict_5_3; // @[LoadQueue.scala 152:68:@15351.4]
  wire  _T_14880; // @[LoadQueue.scala 151:92:@15353.4]
  wire  _T_14881; // @[LoadQueue.scala 152:41:@15354.4]
  wire  _T_14882; // @[LoadQueue.scala 153:30:@15355.4]
  wire  conflict_5_4; // @[LoadQueue.scala 152:68:@15356.4]
  wire  _T_14884; // @[LoadQueue.scala 151:92:@15358.4]
  wire  _T_14885; // @[LoadQueue.scala 152:41:@15359.4]
  wire  _T_14886; // @[LoadQueue.scala 153:30:@15360.4]
  wire  conflict_5_5; // @[LoadQueue.scala 152:68:@15361.4]
  wire  _T_14888; // @[LoadQueue.scala 151:92:@15363.4]
  wire  _T_14889; // @[LoadQueue.scala 152:41:@15364.4]
  wire  _T_14890; // @[LoadQueue.scala 153:30:@15365.4]
  wire  conflict_5_6; // @[LoadQueue.scala 152:68:@15366.4]
  wire  _T_14892; // @[LoadQueue.scala 151:92:@15368.4]
  wire  _T_14893; // @[LoadQueue.scala 152:41:@15369.4]
  wire  _T_14894; // @[LoadQueue.scala 153:30:@15370.4]
  wire  conflict_5_7; // @[LoadQueue.scala 152:68:@15371.4]
  wire  _T_14896; // @[LoadQueue.scala 151:92:@15373.4]
  wire  _T_14897; // @[LoadQueue.scala 152:41:@15374.4]
  wire  _T_14898; // @[LoadQueue.scala 153:30:@15375.4]
  wire  conflict_5_8; // @[LoadQueue.scala 152:68:@15376.4]
  wire  _T_14900; // @[LoadQueue.scala 151:92:@15378.4]
  wire  _T_14901; // @[LoadQueue.scala 152:41:@15379.4]
  wire  _T_14902; // @[LoadQueue.scala 153:30:@15380.4]
  wire  conflict_5_9; // @[LoadQueue.scala 152:68:@15381.4]
  wire  _T_14904; // @[LoadQueue.scala 151:92:@15383.4]
  wire  _T_14905; // @[LoadQueue.scala 152:41:@15384.4]
  wire  _T_14906; // @[LoadQueue.scala 153:30:@15385.4]
  wire  conflict_5_10; // @[LoadQueue.scala 152:68:@15386.4]
  wire  _T_14908; // @[LoadQueue.scala 151:92:@15388.4]
  wire  _T_14909; // @[LoadQueue.scala 152:41:@15389.4]
  wire  _T_14910; // @[LoadQueue.scala 153:30:@15390.4]
  wire  conflict_5_11; // @[LoadQueue.scala 152:68:@15391.4]
  wire  _T_14912; // @[LoadQueue.scala 151:92:@15393.4]
  wire  _T_14913; // @[LoadQueue.scala 152:41:@15394.4]
  wire  _T_14914; // @[LoadQueue.scala 153:30:@15395.4]
  wire  conflict_5_12; // @[LoadQueue.scala 152:68:@15396.4]
  wire  _T_14916; // @[LoadQueue.scala 151:92:@15398.4]
  wire  _T_14917; // @[LoadQueue.scala 152:41:@15399.4]
  wire  _T_14918; // @[LoadQueue.scala 153:30:@15400.4]
  wire  conflict_5_13; // @[LoadQueue.scala 152:68:@15401.4]
  wire  _T_14920; // @[LoadQueue.scala 151:92:@15403.4]
  wire  _T_14921; // @[LoadQueue.scala 152:41:@15404.4]
  wire  _T_14922; // @[LoadQueue.scala 153:30:@15405.4]
  wire  conflict_5_14; // @[LoadQueue.scala 152:68:@15406.4]
  wire  _T_14924; // @[LoadQueue.scala 151:92:@15408.4]
  wire  _T_14925; // @[LoadQueue.scala 152:41:@15409.4]
  wire  _T_14926; // @[LoadQueue.scala 153:30:@15410.4]
  wire  conflict_5_15; // @[LoadQueue.scala 152:68:@15411.4]
  wire  _T_14928; // @[LoadQueue.scala 151:92:@15413.4]
  wire  _T_14929; // @[LoadQueue.scala 152:41:@15414.4]
  wire  _T_14930; // @[LoadQueue.scala 153:30:@15415.4]
  wire  conflict_6_0; // @[LoadQueue.scala 152:68:@15416.4]
  wire  _T_14932; // @[LoadQueue.scala 151:92:@15418.4]
  wire  _T_14933; // @[LoadQueue.scala 152:41:@15419.4]
  wire  _T_14934; // @[LoadQueue.scala 153:30:@15420.4]
  wire  conflict_6_1; // @[LoadQueue.scala 152:68:@15421.4]
  wire  _T_14936; // @[LoadQueue.scala 151:92:@15423.4]
  wire  _T_14937; // @[LoadQueue.scala 152:41:@15424.4]
  wire  _T_14938; // @[LoadQueue.scala 153:30:@15425.4]
  wire  conflict_6_2; // @[LoadQueue.scala 152:68:@15426.4]
  wire  _T_14940; // @[LoadQueue.scala 151:92:@15428.4]
  wire  _T_14941; // @[LoadQueue.scala 152:41:@15429.4]
  wire  _T_14942; // @[LoadQueue.scala 153:30:@15430.4]
  wire  conflict_6_3; // @[LoadQueue.scala 152:68:@15431.4]
  wire  _T_14944; // @[LoadQueue.scala 151:92:@15433.4]
  wire  _T_14945; // @[LoadQueue.scala 152:41:@15434.4]
  wire  _T_14946; // @[LoadQueue.scala 153:30:@15435.4]
  wire  conflict_6_4; // @[LoadQueue.scala 152:68:@15436.4]
  wire  _T_14948; // @[LoadQueue.scala 151:92:@15438.4]
  wire  _T_14949; // @[LoadQueue.scala 152:41:@15439.4]
  wire  _T_14950; // @[LoadQueue.scala 153:30:@15440.4]
  wire  conflict_6_5; // @[LoadQueue.scala 152:68:@15441.4]
  wire  _T_14952; // @[LoadQueue.scala 151:92:@15443.4]
  wire  _T_14953; // @[LoadQueue.scala 152:41:@15444.4]
  wire  _T_14954; // @[LoadQueue.scala 153:30:@15445.4]
  wire  conflict_6_6; // @[LoadQueue.scala 152:68:@15446.4]
  wire  _T_14956; // @[LoadQueue.scala 151:92:@15448.4]
  wire  _T_14957; // @[LoadQueue.scala 152:41:@15449.4]
  wire  _T_14958; // @[LoadQueue.scala 153:30:@15450.4]
  wire  conflict_6_7; // @[LoadQueue.scala 152:68:@15451.4]
  wire  _T_14960; // @[LoadQueue.scala 151:92:@15453.4]
  wire  _T_14961; // @[LoadQueue.scala 152:41:@15454.4]
  wire  _T_14962; // @[LoadQueue.scala 153:30:@15455.4]
  wire  conflict_6_8; // @[LoadQueue.scala 152:68:@15456.4]
  wire  _T_14964; // @[LoadQueue.scala 151:92:@15458.4]
  wire  _T_14965; // @[LoadQueue.scala 152:41:@15459.4]
  wire  _T_14966; // @[LoadQueue.scala 153:30:@15460.4]
  wire  conflict_6_9; // @[LoadQueue.scala 152:68:@15461.4]
  wire  _T_14968; // @[LoadQueue.scala 151:92:@15463.4]
  wire  _T_14969; // @[LoadQueue.scala 152:41:@15464.4]
  wire  _T_14970; // @[LoadQueue.scala 153:30:@15465.4]
  wire  conflict_6_10; // @[LoadQueue.scala 152:68:@15466.4]
  wire  _T_14972; // @[LoadQueue.scala 151:92:@15468.4]
  wire  _T_14973; // @[LoadQueue.scala 152:41:@15469.4]
  wire  _T_14974; // @[LoadQueue.scala 153:30:@15470.4]
  wire  conflict_6_11; // @[LoadQueue.scala 152:68:@15471.4]
  wire  _T_14976; // @[LoadQueue.scala 151:92:@15473.4]
  wire  _T_14977; // @[LoadQueue.scala 152:41:@15474.4]
  wire  _T_14978; // @[LoadQueue.scala 153:30:@15475.4]
  wire  conflict_6_12; // @[LoadQueue.scala 152:68:@15476.4]
  wire  _T_14980; // @[LoadQueue.scala 151:92:@15478.4]
  wire  _T_14981; // @[LoadQueue.scala 152:41:@15479.4]
  wire  _T_14982; // @[LoadQueue.scala 153:30:@15480.4]
  wire  conflict_6_13; // @[LoadQueue.scala 152:68:@15481.4]
  wire  _T_14984; // @[LoadQueue.scala 151:92:@15483.4]
  wire  _T_14985; // @[LoadQueue.scala 152:41:@15484.4]
  wire  _T_14986; // @[LoadQueue.scala 153:30:@15485.4]
  wire  conflict_6_14; // @[LoadQueue.scala 152:68:@15486.4]
  wire  _T_14988; // @[LoadQueue.scala 151:92:@15488.4]
  wire  _T_14989; // @[LoadQueue.scala 152:41:@15489.4]
  wire  _T_14990; // @[LoadQueue.scala 153:30:@15490.4]
  wire  conflict_6_15; // @[LoadQueue.scala 152:68:@15491.4]
  wire  _T_14992; // @[LoadQueue.scala 151:92:@15493.4]
  wire  _T_14993; // @[LoadQueue.scala 152:41:@15494.4]
  wire  _T_14994; // @[LoadQueue.scala 153:30:@15495.4]
  wire  conflict_7_0; // @[LoadQueue.scala 152:68:@15496.4]
  wire  _T_14996; // @[LoadQueue.scala 151:92:@15498.4]
  wire  _T_14997; // @[LoadQueue.scala 152:41:@15499.4]
  wire  _T_14998; // @[LoadQueue.scala 153:30:@15500.4]
  wire  conflict_7_1; // @[LoadQueue.scala 152:68:@15501.4]
  wire  _T_15000; // @[LoadQueue.scala 151:92:@15503.4]
  wire  _T_15001; // @[LoadQueue.scala 152:41:@15504.4]
  wire  _T_15002; // @[LoadQueue.scala 153:30:@15505.4]
  wire  conflict_7_2; // @[LoadQueue.scala 152:68:@15506.4]
  wire  _T_15004; // @[LoadQueue.scala 151:92:@15508.4]
  wire  _T_15005; // @[LoadQueue.scala 152:41:@15509.4]
  wire  _T_15006; // @[LoadQueue.scala 153:30:@15510.4]
  wire  conflict_7_3; // @[LoadQueue.scala 152:68:@15511.4]
  wire  _T_15008; // @[LoadQueue.scala 151:92:@15513.4]
  wire  _T_15009; // @[LoadQueue.scala 152:41:@15514.4]
  wire  _T_15010; // @[LoadQueue.scala 153:30:@15515.4]
  wire  conflict_7_4; // @[LoadQueue.scala 152:68:@15516.4]
  wire  _T_15012; // @[LoadQueue.scala 151:92:@15518.4]
  wire  _T_15013; // @[LoadQueue.scala 152:41:@15519.4]
  wire  _T_15014; // @[LoadQueue.scala 153:30:@15520.4]
  wire  conflict_7_5; // @[LoadQueue.scala 152:68:@15521.4]
  wire  _T_15016; // @[LoadQueue.scala 151:92:@15523.4]
  wire  _T_15017; // @[LoadQueue.scala 152:41:@15524.4]
  wire  _T_15018; // @[LoadQueue.scala 153:30:@15525.4]
  wire  conflict_7_6; // @[LoadQueue.scala 152:68:@15526.4]
  wire  _T_15020; // @[LoadQueue.scala 151:92:@15528.4]
  wire  _T_15021; // @[LoadQueue.scala 152:41:@15529.4]
  wire  _T_15022; // @[LoadQueue.scala 153:30:@15530.4]
  wire  conflict_7_7; // @[LoadQueue.scala 152:68:@15531.4]
  wire  _T_15024; // @[LoadQueue.scala 151:92:@15533.4]
  wire  _T_15025; // @[LoadQueue.scala 152:41:@15534.4]
  wire  _T_15026; // @[LoadQueue.scala 153:30:@15535.4]
  wire  conflict_7_8; // @[LoadQueue.scala 152:68:@15536.4]
  wire  _T_15028; // @[LoadQueue.scala 151:92:@15538.4]
  wire  _T_15029; // @[LoadQueue.scala 152:41:@15539.4]
  wire  _T_15030; // @[LoadQueue.scala 153:30:@15540.4]
  wire  conflict_7_9; // @[LoadQueue.scala 152:68:@15541.4]
  wire  _T_15032; // @[LoadQueue.scala 151:92:@15543.4]
  wire  _T_15033; // @[LoadQueue.scala 152:41:@15544.4]
  wire  _T_15034; // @[LoadQueue.scala 153:30:@15545.4]
  wire  conflict_7_10; // @[LoadQueue.scala 152:68:@15546.4]
  wire  _T_15036; // @[LoadQueue.scala 151:92:@15548.4]
  wire  _T_15037; // @[LoadQueue.scala 152:41:@15549.4]
  wire  _T_15038; // @[LoadQueue.scala 153:30:@15550.4]
  wire  conflict_7_11; // @[LoadQueue.scala 152:68:@15551.4]
  wire  _T_15040; // @[LoadQueue.scala 151:92:@15553.4]
  wire  _T_15041; // @[LoadQueue.scala 152:41:@15554.4]
  wire  _T_15042; // @[LoadQueue.scala 153:30:@15555.4]
  wire  conflict_7_12; // @[LoadQueue.scala 152:68:@15556.4]
  wire  _T_15044; // @[LoadQueue.scala 151:92:@15558.4]
  wire  _T_15045; // @[LoadQueue.scala 152:41:@15559.4]
  wire  _T_15046; // @[LoadQueue.scala 153:30:@15560.4]
  wire  conflict_7_13; // @[LoadQueue.scala 152:68:@15561.4]
  wire  _T_15048; // @[LoadQueue.scala 151:92:@15563.4]
  wire  _T_15049; // @[LoadQueue.scala 152:41:@15564.4]
  wire  _T_15050; // @[LoadQueue.scala 153:30:@15565.4]
  wire  conflict_7_14; // @[LoadQueue.scala 152:68:@15566.4]
  wire  _T_15052; // @[LoadQueue.scala 151:92:@15568.4]
  wire  _T_15053; // @[LoadQueue.scala 152:41:@15569.4]
  wire  _T_15054; // @[LoadQueue.scala 153:30:@15570.4]
  wire  conflict_7_15; // @[LoadQueue.scala 152:68:@15571.4]
  wire  _T_15056; // @[LoadQueue.scala 151:92:@15573.4]
  wire  _T_15057; // @[LoadQueue.scala 152:41:@15574.4]
  wire  _T_15058; // @[LoadQueue.scala 153:30:@15575.4]
  wire  conflict_8_0; // @[LoadQueue.scala 152:68:@15576.4]
  wire  _T_15060; // @[LoadQueue.scala 151:92:@15578.4]
  wire  _T_15061; // @[LoadQueue.scala 152:41:@15579.4]
  wire  _T_15062; // @[LoadQueue.scala 153:30:@15580.4]
  wire  conflict_8_1; // @[LoadQueue.scala 152:68:@15581.4]
  wire  _T_15064; // @[LoadQueue.scala 151:92:@15583.4]
  wire  _T_15065; // @[LoadQueue.scala 152:41:@15584.4]
  wire  _T_15066; // @[LoadQueue.scala 153:30:@15585.4]
  wire  conflict_8_2; // @[LoadQueue.scala 152:68:@15586.4]
  wire  _T_15068; // @[LoadQueue.scala 151:92:@15588.4]
  wire  _T_15069; // @[LoadQueue.scala 152:41:@15589.4]
  wire  _T_15070; // @[LoadQueue.scala 153:30:@15590.4]
  wire  conflict_8_3; // @[LoadQueue.scala 152:68:@15591.4]
  wire  _T_15072; // @[LoadQueue.scala 151:92:@15593.4]
  wire  _T_15073; // @[LoadQueue.scala 152:41:@15594.4]
  wire  _T_15074; // @[LoadQueue.scala 153:30:@15595.4]
  wire  conflict_8_4; // @[LoadQueue.scala 152:68:@15596.4]
  wire  _T_15076; // @[LoadQueue.scala 151:92:@15598.4]
  wire  _T_15077; // @[LoadQueue.scala 152:41:@15599.4]
  wire  _T_15078; // @[LoadQueue.scala 153:30:@15600.4]
  wire  conflict_8_5; // @[LoadQueue.scala 152:68:@15601.4]
  wire  _T_15080; // @[LoadQueue.scala 151:92:@15603.4]
  wire  _T_15081; // @[LoadQueue.scala 152:41:@15604.4]
  wire  _T_15082; // @[LoadQueue.scala 153:30:@15605.4]
  wire  conflict_8_6; // @[LoadQueue.scala 152:68:@15606.4]
  wire  _T_15084; // @[LoadQueue.scala 151:92:@15608.4]
  wire  _T_15085; // @[LoadQueue.scala 152:41:@15609.4]
  wire  _T_15086; // @[LoadQueue.scala 153:30:@15610.4]
  wire  conflict_8_7; // @[LoadQueue.scala 152:68:@15611.4]
  wire  _T_15088; // @[LoadQueue.scala 151:92:@15613.4]
  wire  _T_15089; // @[LoadQueue.scala 152:41:@15614.4]
  wire  _T_15090; // @[LoadQueue.scala 153:30:@15615.4]
  wire  conflict_8_8; // @[LoadQueue.scala 152:68:@15616.4]
  wire  _T_15092; // @[LoadQueue.scala 151:92:@15618.4]
  wire  _T_15093; // @[LoadQueue.scala 152:41:@15619.4]
  wire  _T_15094; // @[LoadQueue.scala 153:30:@15620.4]
  wire  conflict_8_9; // @[LoadQueue.scala 152:68:@15621.4]
  wire  _T_15096; // @[LoadQueue.scala 151:92:@15623.4]
  wire  _T_15097; // @[LoadQueue.scala 152:41:@15624.4]
  wire  _T_15098; // @[LoadQueue.scala 153:30:@15625.4]
  wire  conflict_8_10; // @[LoadQueue.scala 152:68:@15626.4]
  wire  _T_15100; // @[LoadQueue.scala 151:92:@15628.4]
  wire  _T_15101; // @[LoadQueue.scala 152:41:@15629.4]
  wire  _T_15102; // @[LoadQueue.scala 153:30:@15630.4]
  wire  conflict_8_11; // @[LoadQueue.scala 152:68:@15631.4]
  wire  _T_15104; // @[LoadQueue.scala 151:92:@15633.4]
  wire  _T_15105; // @[LoadQueue.scala 152:41:@15634.4]
  wire  _T_15106; // @[LoadQueue.scala 153:30:@15635.4]
  wire  conflict_8_12; // @[LoadQueue.scala 152:68:@15636.4]
  wire  _T_15108; // @[LoadQueue.scala 151:92:@15638.4]
  wire  _T_15109; // @[LoadQueue.scala 152:41:@15639.4]
  wire  _T_15110; // @[LoadQueue.scala 153:30:@15640.4]
  wire  conflict_8_13; // @[LoadQueue.scala 152:68:@15641.4]
  wire  _T_15112; // @[LoadQueue.scala 151:92:@15643.4]
  wire  _T_15113; // @[LoadQueue.scala 152:41:@15644.4]
  wire  _T_15114; // @[LoadQueue.scala 153:30:@15645.4]
  wire  conflict_8_14; // @[LoadQueue.scala 152:68:@15646.4]
  wire  _T_15116; // @[LoadQueue.scala 151:92:@15648.4]
  wire  _T_15117; // @[LoadQueue.scala 152:41:@15649.4]
  wire  _T_15118; // @[LoadQueue.scala 153:30:@15650.4]
  wire  conflict_8_15; // @[LoadQueue.scala 152:68:@15651.4]
  wire  _T_15120; // @[LoadQueue.scala 151:92:@15653.4]
  wire  _T_15121; // @[LoadQueue.scala 152:41:@15654.4]
  wire  _T_15122; // @[LoadQueue.scala 153:30:@15655.4]
  wire  conflict_9_0; // @[LoadQueue.scala 152:68:@15656.4]
  wire  _T_15124; // @[LoadQueue.scala 151:92:@15658.4]
  wire  _T_15125; // @[LoadQueue.scala 152:41:@15659.4]
  wire  _T_15126; // @[LoadQueue.scala 153:30:@15660.4]
  wire  conflict_9_1; // @[LoadQueue.scala 152:68:@15661.4]
  wire  _T_15128; // @[LoadQueue.scala 151:92:@15663.4]
  wire  _T_15129; // @[LoadQueue.scala 152:41:@15664.4]
  wire  _T_15130; // @[LoadQueue.scala 153:30:@15665.4]
  wire  conflict_9_2; // @[LoadQueue.scala 152:68:@15666.4]
  wire  _T_15132; // @[LoadQueue.scala 151:92:@15668.4]
  wire  _T_15133; // @[LoadQueue.scala 152:41:@15669.4]
  wire  _T_15134; // @[LoadQueue.scala 153:30:@15670.4]
  wire  conflict_9_3; // @[LoadQueue.scala 152:68:@15671.4]
  wire  _T_15136; // @[LoadQueue.scala 151:92:@15673.4]
  wire  _T_15137; // @[LoadQueue.scala 152:41:@15674.4]
  wire  _T_15138; // @[LoadQueue.scala 153:30:@15675.4]
  wire  conflict_9_4; // @[LoadQueue.scala 152:68:@15676.4]
  wire  _T_15140; // @[LoadQueue.scala 151:92:@15678.4]
  wire  _T_15141; // @[LoadQueue.scala 152:41:@15679.4]
  wire  _T_15142; // @[LoadQueue.scala 153:30:@15680.4]
  wire  conflict_9_5; // @[LoadQueue.scala 152:68:@15681.4]
  wire  _T_15144; // @[LoadQueue.scala 151:92:@15683.4]
  wire  _T_15145; // @[LoadQueue.scala 152:41:@15684.4]
  wire  _T_15146; // @[LoadQueue.scala 153:30:@15685.4]
  wire  conflict_9_6; // @[LoadQueue.scala 152:68:@15686.4]
  wire  _T_15148; // @[LoadQueue.scala 151:92:@15688.4]
  wire  _T_15149; // @[LoadQueue.scala 152:41:@15689.4]
  wire  _T_15150; // @[LoadQueue.scala 153:30:@15690.4]
  wire  conflict_9_7; // @[LoadQueue.scala 152:68:@15691.4]
  wire  _T_15152; // @[LoadQueue.scala 151:92:@15693.4]
  wire  _T_15153; // @[LoadQueue.scala 152:41:@15694.4]
  wire  _T_15154; // @[LoadQueue.scala 153:30:@15695.4]
  wire  conflict_9_8; // @[LoadQueue.scala 152:68:@15696.4]
  wire  _T_15156; // @[LoadQueue.scala 151:92:@15698.4]
  wire  _T_15157; // @[LoadQueue.scala 152:41:@15699.4]
  wire  _T_15158; // @[LoadQueue.scala 153:30:@15700.4]
  wire  conflict_9_9; // @[LoadQueue.scala 152:68:@15701.4]
  wire  _T_15160; // @[LoadQueue.scala 151:92:@15703.4]
  wire  _T_15161; // @[LoadQueue.scala 152:41:@15704.4]
  wire  _T_15162; // @[LoadQueue.scala 153:30:@15705.4]
  wire  conflict_9_10; // @[LoadQueue.scala 152:68:@15706.4]
  wire  _T_15164; // @[LoadQueue.scala 151:92:@15708.4]
  wire  _T_15165; // @[LoadQueue.scala 152:41:@15709.4]
  wire  _T_15166; // @[LoadQueue.scala 153:30:@15710.4]
  wire  conflict_9_11; // @[LoadQueue.scala 152:68:@15711.4]
  wire  _T_15168; // @[LoadQueue.scala 151:92:@15713.4]
  wire  _T_15169; // @[LoadQueue.scala 152:41:@15714.4]
  wire  _T_15170; // @[LoadQueue.scala 153:30:@15715.4]
  wire  conflict_9_12; // @[LoadQueue.scala 152:68:@15716.4]
  wire  _T_15172; // @[LoadQueue.scala 151:92:@15718.4]
  wire  _T_15173; // @[LoadQueue.scala 152:41:@15719.4]
  wire  _T_15174; // @[LoadQueue.scala 153:30:@15720.4]
  wire  conflict_9_13; // @[LoadQueue.scala 152:68:@15721.4]
  wire  _T_15176; // @[LoadQueue.scala 151:92:@15723.4]
  wire  _T_15177; // @[LoadQueue.scala 152:41:@15724.4]
  wire  _T_15178; // @[LoadQueue.scala 153:30:@15725.4]
  wire  conflict_9_14; // @[LoadQueue.scala 152:68:@15726.4]
  wire  _T_15180; // @[LoadQueue.scala 151:92:@15728.4]
  wire  _T_15181; // @[LoadQueue.scala 152:41:@15729.4]
  wire  _T_15182; // @[LoadQueue.scala 153:30:@15730.4]
  wire  conflict_9_15; // @[LoadQueue.scala 152:68:@15731.4]
  wire  _T_15184; // @[LoadQueue.scala 151:92:@15733.4]
  wire  _T_15185; // @[LoadQueue.scala 152:41:@15734.4]
  wire  _T_15186; // @[LoadQueue.scala 153:30:@15735.4]
  wire  conflict_10_0; // @[LoadQueue.scala 152:68:@15736.4]
  wire  _T_15188; // @[LoadQueue.scala 151:92:@15738.4]
  wire  _T_15189; // @[LoadQueue.scala 152:41:@15739.4]
  wire  _T_15190; // @[LoadQueue.scala 153:30:@15740.4]
  wire  conflict_10_1; // @[LoadQueue.scala 152:68:@15741.4]
  wire  _T_15192; // @[LoadQueue.scala 151:92:@15743.4]
  wire  _T_15193; // @[LoadQueue.scala 152:41:@15744.4]
  wire  _T_15194; // @[LoadQueue.scala 153:30:@15745.4]
  wire  conflict_10_2; // @[LoadQueue.scala 152:68:@15746.4]
  wire  _T_15196; // @[LoadQueue.scala 151:92:@15748.4]
  wire  _T_15197; // @[LoadQueue.scala 152:41:@15749.4]
  wire  _T_15198; // @[LoadQueue.scala 153:30:@15750.4]
  wire  conflict_10_3; // @[LoadQueue.scala 152:68:@15751.4]
  wire  _T_15200; // @[LoadQueue.scala 151:92:@15753.4]
  wire  _T_15201; // @[LoadQueue.scala 152:41:@15754.4]
  wire  _T_15202; // @[LoadQueue.scala 153:30:@15755.4]
  wire  conflict_10_4; // @[LoadQueue.scala 152:68:@15756.4]
  wire  _T_15204; // @[LoadQueue.scala 151:92:@15758.4]
  wire  _T_15205; // @[LoadQueue.scala 152:41:@15759.4]
  wire  _T_15206; // @[LoadQueue.scala 153:30:@15760.4]
  wire  conflict_10_5; // @[LoadQueue.scala 152:68:@15761.4]
  wire  _T_15208; // @[LoadQueue.scala 151:92:@15763.4]
  wire  _T_15209; // @[LoadQueue.scala 152:41:@15764.4]
  wire  _T_15210; // @[LoadQueue.scala 153:30:@15765.4]
  wire  conflict_10_6; // @[LoadQueue.scala 152:68:@15766.4]
  wire  _T_15212; // @[LoadQueue.scala 151:92:@15768.4]
  wire  _T_15213; // @[LoadQueue.scala 152:41:@15769.4]
  wire  _T_15214; // @[LoadQueue.scala 153:30:@15770.4]
  wire  conflict_10_7; // @[LoadQueue.scala 152:68:@15771.4]
  wire  _T_15216; // @[LoadQueue.scala 151:92:@15773.4]
  wire  _T_15217; // @[LoadQueue.scala 152:41:@15774.4]
  wire  _T_15218; // @[LoadQueue.scala 153:30:@15775.4]
  wire  conflict_10_8; // @[LoadQueue.scala 152:68:@15776.4]
  wire  _T_15220; // @[LoadQueue.scala 151:92:@15778.4]
  wire  _T_15221; // @[LoadQueue.scala 152:41:@15779.4]
  wire  _T_15222; // @[LoadQueue.scala 153:30:@15780.4]
  wire  conflict_10_9; // @[LoadQueue.scala 152:68:@15781.4]
  wire  _T_15224; // @[LoadQueue.scala 151:92:@15783.4]
  wire  _T_15225; // @[LoadQueue.scala 152:41:@15784.4]
  wire  _T_15226; // @[LoadQueue.scala 153:30:@15785.4]
  wire  conflict_10_10; // @[LoadQueue.scala 152:68:@15786.4]
  wire  _T_15228; // @[LoadQueue.scala 151:92:@15788.4]
  wire  _T_15229; // @[LoadQueue.scala 152:41:@15789.4]
  wire  _T_15230; // @[LoadQueue.scala 153:30:@15790.4]
  wire  conflict_10_11; // @[LoadQueue.scala 152:68:@15791.4]
  wire  _T_15232; // @[LoadQueue.scala 151:92:@15793.4]
  wire  _T_15233; // @[LoadQueue.scala 152:41:@15794.4]
  wire  _T_15234; // @[LoadQueue.scala 153:30:@15795.4]
  wire  conflict_10_12; // @[LoadQueue.scala 152:68:@15796.4]
  wire  _T_15236; // @[LoadQueue.scala 151:92:@15798.4]
  wire  _T_15237; // @[LoadQueue.scala 152:41:@15799.4]
  wire  _T_15238; // @[LoadQueue.scala 153:30:@15800.4]
  wire  conflict_10_13; // @[LoadQueue.scala 152:68:@15801.4]
  wire  _T_15240; // @[LoadQueue.scala 151:92:@15803.4]
  wire  _T_15241; // @[LoadQueue.scala 152:41:@15804.4]
  wire  _T_15242; // @[LoadQueue.scala 153:30:@15805.4]
  wire  conflict_10_14; // @[LoadQueue.scala 152:68:@15806.4]
  wire  _T_15244; // @[LoadQueue.scala 151:92:@15808.4]
  wire  _T_15245; // @[LoadQueue.scala 152:41:@15809.4]
  wire  _T_15246; // @[LoadQueue.scala 153:30:@15810.4]
  wire  conflict_10_15; // @[LoadQueue.scala 152:68:@15811.4]
  wire  _T_15248; // @[LoadQueue.scala 151:92:@15813.4]
  wire  _T_15249; // @[LoadQueue.scala 152:41:@15814.4]
  wire  _T_15250; // @[LoadQueue.scala 153:30:@15815.4]
  wire  conflict_11_0; // @[LoadQueue.scala 152:68:@15816.4]
  wire  _T_15252; // @[LoadQueue.scala 151:92:@15818.4]
  wire  _T_15253; // @[LoadQueue.scala 152:41:@15819.4]
  wire  _T_15254; // @[LoadQueue.scala 153:30:@15820.4]
  wire  conflict_11_1; // @[LoadQueue.scala 152:68:@15821.4]
  wire  _T_15256; // @[LoadQueue.scala 151:92:@15823.4]
  wire  _T_15257; // @[LoadQueue.scala 152:41:@15824.4]
  wire  _T_15258; // @[LoadQueue.scala 153:30:@15825.4]
  wire  conflict_11_2; // @[LoadQueue.scala 152:68:@15826.4]
  wire  _T_15260; // @[LoadQueue.scala 151:92:@15828.4]
  wire  _T_15261; // @[LoadQueue.scala 152:41:@15829.4]
  wire  _T_15262; // @[LoadQueue.scala 153:30:@15830.4]
  wire  conflict_11_3; // @[LoadQueue.scala 152:68:@15831.4]
  wire  _T_15264; // @[LoadQueue.scala 151:92:@15833.4]
  wire  _T_15265; // @[LoadQueue.scala 152:41:@15834.4]
  wire  _T_15266; // @[LoadQueue.scala 153:30:@15835.4]
  wire  conflict_11_4; // @[LoadQueue.scala 152:68:@15836.4]
  wire  _T_15268; // @[LoadQueue.scala 151:92:@15838.4]
  wire  _T_15269; // @[LoadQueue.scala 152:41:@15839.4]
  wire  _T_15270; // @[LoadQueue.scala 153:30:@15840.4]
  wire  conflict_11_5; // @[LoadQueue.scala 152:68:@15841.4]
  wire  _T_15272; // @[LoadQueue.scala 151:92:@15843.4]
  wire  _T_15273; // @[LoadQueue.scala 152:41:@15844.4]
  wire  _T_15274; // @[LoadQueue.scala 153:30:@15845.4]
  wire  conflict_11_6; // @[LoadQueue.scala 152:68:@15846.4]
  wire  _T_15276; // @[LoadQueue.scala 151:92:@15848.4]
  wire  _T_15277; // @[LoadQueue.scala 152:41:@15849.4]
  wire  _T_15278; // @[LoadQueue.scala 153:30:@15850.4]
  wire  conflict_11_7; // @[LoadQueue.scala 152:68:@15851.4]
  wire  _T_15280; // @[LoadQueue.scala 151:92:@15853.4]
  wire  _T_15281; // @[LoadQueue.scala 152:41:@15854.4]
  wire  _T_15282; // @[LoadQueue.scala 153:30:@15855.4]
  wire  conflict_11_8; // @[LoadQueue.scala 152:68:@15856.4]
  wire  _T_15284; // @[LoadQueue.scala 151:92:@15858.4]
  wire  _T_15285; // @[LoadQueue.scala 152:41:@15859.4]
  wire  _T_15286; // @[LoadQueue.scala 153:30:@15860.4]
  wire  conflict_11_9; // @[LoadQueue.scala 152:68:@15861.4]
  wire  _T_15288; // @[LoadQueue.scala 151:92:@15863.4]
  wire  _T_15289; // @[LoadQueue.scala 152:41:@15864.4]
  wire  _T_15290; // @[LoadQueue.scala 153:30:@15865.4]
  wire  conflict_11_10; // @[LoadQueue.scala 152:68:@15866.4]
  wire  _T_15292; // @[LoadQueue.scala 151:92:@15868.4]
  wire  _T_15293; // @[LoadQueue.scala 152:41:@15869.4]
  wire  _T_15294; // @[LoadQueue.scala 153:30:@15870.4]
  wire  conflict_11_11; // @[LoadQueue.scala 152:68:@15871.4]
  wire  _T_15296; // @[LoadQueue.scala 151:92:@15873.4]
  wire  _T_15297; // @[LoadQueue.scala 152:41:@15874.4]
  wire  _T_15298; // @[LoadQueue.scala 153:30:@15875.4]
  wire  conflict_11_12; // @[LoadQueue.scala 152:68:@15876.4]
  wire  _T_15300; // @[LoadQueue.scala 151:92:@15878.4]
  wire  _T_15301; // @[LoadQueue.scala 152:41:@15879.4]
  wire  _T_15302; // @[LoadQueue.scala 153:30:@15880.4]
  wire  conflict_11_13; // @[LoadQueue.scala 152:68:@15881.4]
  wire  _T_15304; // @[LoadQueue.scala 151:92:@15883.4]
  wire  _T_15305; // @[LoadQueue.scala 152:41:@15884.4]
  wire  _T_15306; // @[LoadQueue.scala 153:30:@15885.4]
  wire  conflict_11_14; // @[LoadQueue.scala 152:68:@15886.4]
  wire  _T_15308; // @[LoadQueue.scala 151:92:@15888.4]
  wire  _T_15309; // @[LoadQueue.scala 152:41:@15889.4]
  wire  _T_15310; // @[LoadQueue.scala 153:30:@15890.4]
  wire  conflict_11_15; // @[LoadQueue.scala 152:68:@15891.4]
  wire  _T_15312; // @[LoadQueue.scala 151:92:@15893.4]
  wire  _T_15313; // @[LoadQueue.scala 152:41:@15894.4]
  wire  _T_15314; // @[LoadQueue.scala 153:30:@15895.4]
  wire  conflict_12_0; // @[LoadQueue.scala 152:68:@15896.4]
  wire  _T_15316; // @[LoadQueue.scala 151:92:@15898.4]
  wire  _T_15317; // @[LoadQueue.scala 152:41:@15899.4]
  wire  _T_15318; // @[LoadQueue.scala 153:30:@15900.4]
  wire  conflict_12_1; // @[LoadQueue.scala 152:68:@15901.4]
  wire  _T_15320; // @[LoadQueue.scala 151:92:@15903.4]
  wire  _T_15321; // @[LoadQueue.scala 152:41:@15904.4]
  wire  _T_15322; // @[LoadQueue.scala 153:30:@15905.4]
  wire  conflict_12_2; // @[LoadQueue.scala 152:68:@15906.4]
  wire  _T_15324; // @[LoadQueue.scala 151:92:@15908.4]
  wire  _T_15325; // @[LoadQueue.scala 152:41:@15909.4]
  wire  _T_15326; // @[LoadQueue.scala 153:30:@15910.4]
  wire  conflict_12_3; // @[LoadQueue.scala 152:68:@15911.4]
  wire  _T_15328; // @[LoadQueue.scala 151:92:@15913.4]
  wire  _T_15329; // @[LoadQueue.scala 152:41:@15914.4]
  wire  _T_15330; // @[LoadQueue.scala 153:30:@15915.4]
  wire  conflict_12_4; // @[LoadQueue.scala 152:68:@15916.4]
  wire  _T_15332; // @[LoadQueue.scala 151:92:@15918.4]
  wire  _T_15333; // @[LoadQueue.scala 152:41:@15919.4]
  wire  _T_15334; // @[LoadQueue.scala 153:30:@15920.4]
  wire  conflict_12_5; // @[LoadQueue.scala 152:68:@15921.4]
  wire  _T_15336; // @[LoadQueue.scala 151:92:@15923.4]
  wire  _T_15337; // @[LoadQueue.scala 152:41:@15924.4]
  wire  _T_15338; // @[LoadQueue.scala 153:30:@15925.4]
  wire  conflict_12_6; // @[LoadQueue.scala 152:68:@15926.4]
  wire  _T_15340; // @[LoadQueue.scala 151:92:@15928.4]
  wire  _T_15341; // @[LoadQueue.scala 152:41:@15929.4]
  wire  _T_15342; // @[LoadQueue.scala 153:30:@15930.4]
  wire  conflict_12_7; // @[LoadQueue.scala 152:68:@15931.4]
  wire  _T_15344; // @[LoadQueue.scala 151:92:@15933.4]
  wire  _T_15345; // @[LoadQueue.scala 152:41:@15934.4]
  wire  _T_15346; // @[LoadQueue.scala 153:30:@15935.4]
  wire  conflict_12_8; // @[LoadQueue.scala 152:68:@15936.4]
  wire  _T_15348; // @[LoadQueue.scala 151:92:@15938.4]
  wire  _T_15349; // @[LoadQueue.scala 152:41:@15939.4]
  wire  _T_15350; // @[LoadQueue.scala 153:30:@15940.4]
  wire  conflict_12_9; // @[LoadQueue.scala 152:68:@15941.4]
  wire  _T_15352; // @[LoadQueue.scala 151:92:@15943.4]
  wire  _T_15353; // @[LoadQueue.scala 152:41:@15944.4]
  wire  _T_15354; // @[LoadQueue.scala 153:30:@15945.4]
  wire  conflict_12_10; // @[LoadQueue.scala 152:68:@15946.4]
  wire  _T_15356; // @[LoadQueue.scala 151:92:@15948.4]
  wire  _T_15357; // @[LoadQueue.scala 152:41:@15949.4]
  wire  _T_15358; // @[LoadQueue.scala 153:30:@15950.4]
  wire  conflict_12_11; // @[LoadQueue.scala 152:68:@15951.4]
  wire  _T_15360; // @[LoadQueue.scala 151:92:@15953.4]
  wire  _T_15361; // @[LoadQueue.scala 152:41:@15954.4]
  wire  _T_15362; // @[LoadQueue.scala 153:30:@15955.4]
  wire  conflict_12_12; // @[LoadQueue.scala 152:68:@15956.4]
  wire  _T_15364; // @[LoadQueue.scala 151:92:@15958.4]
  wire  _T_15365; // @[LoadQueue.scala 152:41:@15959.4]
  wire  _T_15366; // @[LoadQueue.scala 153:30:@15960.4]
  wire  conflict_12_13; // @[LoadQueue.scala 152:68:@15961.4]
  wire  _T_15368; // @[LoadQueue.scala 151:92:@15963.4]
  wire  _T_15369; // @[LoadQueue.scala 152:41:@15964.4]
  wire  _T_15370; // @[LoadQueue.scala 153:30:@15965.4]
  wire  conflict_12_14; // @[LoadQueue.scala 152:68:@15966.4]
  wire  _T_15372; // @[LoadQueue.scala 151:92:@15968.4]
  wire  _T_15373; // @[LoadQueue.scala 152:41:@15969.4]
  wire  _T_15374; // @[LoadQueue.scala 153:30:@15970.4]
  wire  conflict_12_15; // @[LoadQueue.scala 152:68:@15971.4]
  wire  _T_15376; // @[LoadQueue.scala 151:92:@15973.4]
  wire  _T_15377; // @[LoadQueue.scala 152:41:@15974.4]
  wire  _T_15378; // @[LoadQueue.scala 153:30:@15975.4]
  wire  conflict_13_0; // @[LoadQueue.scala 152:68:@15976.4]
  wire  _T_15380; // @[LoadQueue.scala 151:92:@15978.4]
  wire  _T_15381; // @[LoadQueue.scala 152:41:@15979.4]
  wire  _T_15382; // @[LoadQueue.scala 153:30:@15980.4]
  wire  conflict_13_1; // @[LoadQueue.scala 152:68:@15981.4]
  wire  _T_15384; // @[LoadQueue.scala 151:92:@15983.4]
  wire  _T_15385; // @[LoadQueue.scala 152:41:@15984.4]
  wire  _T_15386; // @[LoadQueue.scala 153:30:@15985.4]
  wire  conflict_13_2; // @[LoadQueue.scala 152:68:@15986.4]
  wire  _T_15388; // @[LoadQueue.scala 151:92:@15988.4]
  wire  _T_15389; // @[LoadQueue.scala 152:41:@15989.4]
  wire  _T_15390; // @[LoadQueue.scala 153:30:@15990.4]
  wire  conflict_13_3; // @[LoadQueue.scala 152:68:@15991.4]
  wire  _T_15392; // @[LoadQueue.scala 151:92:@15993.4]
  wire  _T_15393; // @[LoadQueue.scala 152:41:@15994.4]
  wire  _T_15394; // @[LoadQueue.scala 153:30:@15995.4]
  wire  conflict_13_4; // @[LoadQueue.scala 152:68:@15996.4]
  wire  _T_15396; // @[LoadQueue.scala 151:92:@15998.4]
  wire  _T_15397; // @[LoadQueue.scala 152:41:@15999.4]
  wire  _T_15398; // @[LoadQueue.scala 153:30:@16000.4]
  wire  conflict_13_5; // @[LoadQueue.scala 152:68:@16001.4]
  wire  _T_15400; // @[LoadQueue.scala 151:92:@16003.4]
  wire  _T_15401; // @[LoadQueue.scala 152:41:@16004.4]
  wire  _T_15402; // @[LoadQueue.scala 153:30:@16005.4]
  wire  conflict_13_6; // @[LoadQueue.scala 152:68:@16006.4]
  wire  _T_15404; // @[LoadQueue.scala 151:92:@16008.4]
  wire  _T_15405; // @[LoadQueue.scala 152:41:@16009.4]
  wire  _T_15406; // @[LoadQueue.scala 153:30:@16010.4]
  wire  conflict_13_7; // @[LoadQueue.scala 152:68:@16011.4]
  wire  _T_15408; // @[LoadQueue.scala 151:92:@16013.4]
  wire  _T_15409; // @[LoadQueue.scala 152:41:@16014.4]
  wire  _T_15410; // @[LoadQueue.scala 153:30:@16015.4]
  wire  conflict_13_8; // @[LoadQueue.scala 152:68:@16016.4]
  wire  _T_15412; // @[LoadQueue.scala 151:92:@16018.4]
  wire  _T_15413; // @[LoadQueue.scala 152:41:@16019.4]
  wire  _T_15414; // @[LoadQueue.scala 153:30:@16020.4]
  wire  conflict_13_9; // @[LoadQueue.scala 152:68:@16021.4]
  wire  _T_15416; // @[LoadQueue.scala 151:92:@16023.4]
  wire  _T_15417; // @[LoadQueue.scala 152:41:@16024.4]
  wire  _T_15418; // @[LoadQueue.scala 153:30:@16025.4]
  wire  conflict_13_10; // @[LoadQueue.scala 152:68:@16026.4]
  wire  _T_15420; // @[LoadQueue.scala 151:92:@16028.4]
  wire  _T_15421; // @[LoadQueue.scala 152:41:@16029.4]
  wire  _T_15422; // @[LoadQueue.scala 153:30:@16030.4]
  wire  conflict_13_11; // @[LoadQueue.scala 152:68:@16031.4]
  wire  _T_15424; // @[LoadQueue.scala 151:92:@16033.4]
  wire  _T_15425; // @[LoadQueue.scala 152:41:@16034.4]
  wire  _T_15426; // @[LoadQueue.scala 153:30:@16035.4]
  wire  conflict_13_12; // @[LoadQueue.scala 152:68:@16036.4]
  wire  _T_15428; // @[LoadQueue.scala 151:92:@16038.4]
  wire  _T_15429; // @[LoadQueue.scala 152:41:@16039.4]
  wire  _T_15430; // @[LoadQueue.scala 153:30:@16040.4]
  wire  conflict_13_13; // @[LoadQueue.scala 152:68:@16041.4]
  wire  _T_15432; // @[LoadQueue.scala 151:92:@16043.4]
  wire  _T_15433; // @[LoadQueue.scala 152:41:@16044.4]
  wire  _T_15434; // @[LoadQueue.scala 153:30:@16045.4]
  wire  conflict_13_14; // @[LoadQueue.scala 152:68:@16046.4]
  wire  _T_15436; // @[LoadQueue.scala 151:92:@16048.4]
  wire  _T_15437; // @[LoadQueue.scala 152:41:@16049.4]
  wire  _T_15438; // @[LoadQueue.scala 153:30:@16050.4]
  wire  conflict_13_15; // @[LoadQueue.scala 152:68:@16051.4]
  wire  _T_15440; // @[LoadQueue.scala 151:92:@16053.4]
  wire  _T_15441; // @[LoadQueue.scala 152:41:@16054.4]
  wire  _T_15442; // @[LoadQueue.scala 153:30:@16055.4]
  wire  conflict_14_0; // @[LoadQueue.scala 152:68:@16056.4]
  wire  _T_15444; // @[LoadQueue.scala 151:92:@16058.4]
  wire  _T_15445; // @[LoadQueue.scala 152:41:@16059.4]
  wire  _T_15446; // @[LoadQueue.scala 153:30:@16060.4]
  wire  conflict_14_1; // @[LoadQueue.scala 152:68:@16061.4]
  wire  _T_15448; // @[LoadQueue.scala 151:92:@16063.4]
  wire  _T_15449; // @[LoadQueue.scala 152:41:@16064.4]
  wire  _T_15450; // @[LoadQueue.scala 153:30:@16065.4]
  wire  conflict_14_2; // @[LoadQueue.scala 152:68:@16066.4]
  wire  _T_15452; // @[LoadQueue.scala 151:92:@16068.4]
  wire  _T_15453; // @[LoadQueue.scala 152:41:@16069.4]
  wire  _T_15454; // @[LoadQueue.scala 153:30:@16070.4]
  wire  conflict_14_3; // @[LoadQueue.scala 152:68:@16071.4]
  wire  _T_15456; // @[LoadQueue.scala 151:92:@16073.4]
  wire  _T_15457; // @[LoadQueue.scala 152:41:@16074.4]
  wire  _T_15458; // @[LoadQueue.scala 153:30:@16075.4]
  wire  conflict_14_4; // @[LoadQueue.scala 152:68:@16076.4]
  wire  _T_15460; // @[LoadQueue.scala 151:92:@16078.4]
  wire  _T_15461; // @[LoadQueue.scala 152:41:@16079.4]
  wire  _T_15462; // @[LoadQueue.scala 153:30:@16080.4]
  wire  conflict_14_5; // @[LoadQueue.scala 152:68:@16081.4]
  wire  _T_15464; // @[LoadQueue.scala 151:92:@16083.4]
  wire  _T_15465; // @[LoadQueue.scala 152:41:@16084.4]
  wire  _T_15466; // @[LoadQueue.scala 153:30:@16085.4]
  wire  conflict_14_6; // @[LoadQueue.scala 152:68:@16086.4]
  wire  _T_15468; // @[LoadQueue.scala 151:92:@16088.4]
  wire  _T_15469; // @[LoadQueue.scala 152:41:@16089.4]
  wire  _T_15470; // @[LoadQueue.scala 153:30:@16090.4]
  wire  conflict_14_7; // @[LoadQueue.scala 152:68:@16091.4]
  wire  _T_15472; // @[LoadQueue.scala 151:92:@16093.4]
  wire  _T_15473; // @[LoadQueue.scala 152:41:@16094.4]
  wire  _T_15474; // @[LoadQueue.scala 153:30:@16095.4]
  wire  conflict_14_8; // @[LoadQueue.scala 152:68:@16096.4]
  wire  _T_15476; // @[LoadQueue.scala 151:92:@16098.4]
  wire  _T_15477; // @[LoadQueue.scala 152:41:@16099.4]
  wire  _T_15478; // @[LoadQueue.scala 153:30:@16100.4]
  wire  conflict_14_9; // @[LoadQueue.scala 152:68:@16101.4]
  wire  _T_15480; // @[LoadQueue.scala 151:92:@16103.4]
  wire  _T_15481; // @[LoadQueue.scala 152:41:@16104.4]
  wire  _T_15482; // @[LoadQueue.scala 153:30:@16105.4]
  wire  conflict_14_10; // @[LoadQueue.scala 152:68:@16106.4]
  wire  _T_15484; // @[LoadQueue.scala 151:92:@16108.4]
  wire  _T_15485; // @[LoadQueue.scala 152:41:@16109.4]
  wire  _T_15486; // @[LoadQueue.scala 153:30:@16110.4]
  wire  conflict_14_11; // @[LoadQueue.scala 152:68:@16111.4]
  wire  _T_15488; // @[LoadQueue.scala 151:92:@16113.4]
  wire  _T_15489; // @[LoadQueue.scala 152:41:@16114.4]
  wire  _T_15490; // @[LoadQueue.scala 153:30:@16115.4]
  wire  conflict_14_12; // @[LoadQueue.scala 152:68:@16116.4]
  wire  _T_15492; // @[LoadQueue.scala 151:92:@16118.4]
  wire  _T_15493; // @[LoadQueue.scala 152:41:@16119.4]
  wire  _T_15494; // @[LoadQueue.scala 153:30:@16120.4]
  wire  conflict_14_13; // @[LoadQueue.scala 152:68:@16121.4]
  wire  _T_15496; // @[LoadQueue.scala 151:92:@16123.4]
  wire  _T_15497; // @[LoadQueue.scala 152:41:@16124.4]
  wire  _T_15498; // @[LoadQueue.scala 153:30:@16125.4]
  wire  conflict_14_14; // @[LoadQueue.scala 152:68:@16126.4]
  wire  _T_15500; // @[LoadQueue.scala 151:92:@16128.4]
  wire  _T_15501; // @[LoadQueue.scala 152:41:@16129.4]
  wire  _T_15502; // @[LoadQueue.scala 153:30:@16130.4]
  wire  conflict_14_15; // @[LoadQueue.scala 152:68:@16131.4]
  wire  _T_15504; // @[LoadQueue.scala 151:92:@16133.4]
  wire  _T_15505; // @[LoadQueue.scala 152:41:@16134.4]
  wire  _T_15506; // @[LoadQueue.scala 153:30:@16135.4]
  wire  conflict_15_0; // @[LoadQueue.scala 152:68:@16136.4]
  wire  _T_15508; // @[LoadQueue.scala 151:92:@16138.4]
  wire  _T_15509; // @[LoadQueue.scala 152:41:@16139.4]
  wire  _T_15510; // @[LoadQueue.scala 153:30:@16140.4]
  wire  conflict_15_1; // @[LoadQueue.scala 152:68:@16141.4]
  wire  _T_15512; // @[LoadQueue.scala 151:92:@16143.4]
  wire  _T_15513; // @[LoadQueue.scala 152:41:@16144.4]
  wire  _T_15514; // @[LoadQueue.scala 153:30:@16145.4]
  wire  conflict_15_2; // @[LoadQueue.scala 152:68:@16146.4]
  wire  _T_15516; // @[LoadQueue.scala 151:92:@16148.4]
  wire  _T_15517; // @[LoadQueue.scala 152:41:@16149.4]
  wire  _T_15518; // @[LoadQueue.scala 153:30:@16150.4]
  wire  conflict_15_3; // @[LoadQueue.scala 152:68:@16151.4]
  wire  _T_15520; // @[LoadQueue.scala 151:92:@16153.4]
  wire  _T_15521; // @[LoadQueue.scala 152:41:@16154.4]
  wire  _T_15522; // @[LoadQueue.scala 153:30:@16155.4]
  wire  conflict_15_4; // @[LoadQueue.scala 152:68:@16156.4]
  wire  _T_15524; // @[LoadQueue.scala 151:92:@16158.4]
  wire  _T_15525; // @[LoadQueue.scala 152:41:@16159.4]
  wire  _T_15526; // @[LoadQueue.scala 153:30:@16160.4]
  wire  conflict_15_5; // @[LoadQueue.scala 152:68:@16161.4]
  wire  _T_15528; // @[LoadQueue.scala 151:92:@16163.4]
  wire  _T_15529; // @[LoadQueue.scala 152:41:@16164.4]
  wire  _T_15530; // @[LoadQueue.scala 153:30:@16165.4]
  wire  conflict_15_6; // @[LoadQueue.scala 152:68:@16166.4]
  wire  _T_15532; // @[LoadQueue.scala 151:92:@16168.4]
  wire  _T_15533; // @[LoadQueue.scala 152:41:@16169.4]
  wire  _T_15534; // @[LoadQueue.scala 153:30:@16170.4]
  wire  conflict_15_7; // @[LoadQueue.scala 152:68:@16171.4]
  wire  _T_15536; // @[LoadQueue.scala 151:92:@16173.4]
  wire  _T_15537; // @[LoadQueue.scala 152:41:@16174.4]
  wire  _T_15538; // @[LoadQueue.scala 153:30:@16175.4]
  wire  conflict_15_8; // @[LoadQueue.scala 152:68:@16176.4]
  wire  _T_15540; // @[LoadQueue.scala 151:92:@16178.4]
  wire  _T_15541; // @[LoadQueue.scala 152:41:@16179.4]
  wire  _T_15542; // @[LoadQueue.scala 153:30:@16180.4]
  wire  conflict_15_9; // @[LoadQueue.scala 152:68:@16181.4]
  wire  _T_15544; // @[LoadQueue.scala 151:92:@16183.4]
  wire  _T_15545; // @[LoadQueue.scala 152:41:@16184.4]
  wire  _T_15546; // @[LoadQueue.scala 153:30:@16185.4]
  wire  conflict_15_10; // @[LoadQueue.scala 152:68:@16186.4]
  wire  _T_15548; // @[LoadQueue.scala 151:92:@16188.4]
  wire  _T_15549; // @[LoadQueue.scala 152:41:@16189.4]
  wire  _T_15550; // @[LoadQueue.scala 153:30:@16190.4]
  wire  conflict_15_11; // @[LoadQueue.scala 152:68:@16191.4]
  wire  _T_15552; // @[LoadQueue.scala 151:92:@16193.4]
  wire  _T_15553; // @[LoadQueue.scala 152:41:@16194.4]
  wire  _T_15554; // @[LoadQueue.scala 153:30:@16195.4]
  wire  conflict_15_12; // @[LoadQueue.scala 152:68:@16196.4]
  wire  _T_15556; // @[LoadQueue.scala 151:92:@16198.4]
  wire  _T_15557; // @[LoadQueue.scala 152:41:@16199.4]
  wire  _T_15558; // @[LoadQueue.scala 153:30:@16200.4]
  wire  conflict_15_13; // @[LoadQueue.scala 152:68:@16201.4]
  wire  _T_15560; // @[LoadQueue.scala 151:92:@16203.4]
  wire  _T_15561; // @[LoadQueue.scala 152:41:@16204.4]
  wire  _T_15562; // @[LoadQueue.scala 153:30:@16205.4]
  wire  conflict_15_14; // @[LoadQueue.scala 152:68:@16206.4]
  wire  _T_15564; // @[LoadQueue.scala 151:92:@16208.4]
  wire  _T_15565; // @[LoadQueue.scala 152:41:@16209.4]
  wire  _T_15566; // @[LoadQueue.scala 153:30:@16210.4]
  wire  conflict_15_15; // @[LoadQueue.scala 152:68:@16211.4]
  wire  _T_16799; // @[LoadQueue.scala 163:13:@16214.4]
  wire  storeAddrNotKnownFlags_0_0; // @[LoadQueue.scala 163:19:@16215.4]
  wire  _T_16802; // @[LoadQueue.scala 163:13:@16216.4]
  wire  storeAddrNotKnownFlags_0_1; // @[LoadQueue.scala 163:19:@16217.4]
  wire  _T_16805; // @[LoadQueue.scala 163:13:@16218.4]
  wire  storeAddrNotKnownFlags_0_2; // @[LoadQueue.scala 163:19:@16219.4]
  wire  _T_16808; // @[LoadQueue.scala 163:13:@16220.4]
  wire  storeAddrNotKnownFlags_0_3; // @[LoadQueue.scala 163:19:@16221.4]
  wire  _T_16811; // @[LoadQueue.scala 163:13:@16222.4]
  wire  storeAddrNotKnownFlags_0_4; // @[LoadQueue.scala 163:19:@16223.4]
  wire  _T_16814; // @[LoadQueue.scala 163:13:@16224.4]
  wire  storeAddrNotKnownFlags_0_5; // @[LoadQueue.scala 163:19:@16225.4]
  wire  _T_16817; // @[LoadQueue.scala 163:13:@16226.4]
  wire  storeAddrNotKnownFlags_0_6; // @[LoadQueue.scala 163:19:@16227.4]
  wire  _T_16820; // @[LoadQueue.scala 163:13:@16228.4]
  wire  storeAddrNotKnownFlags_0_7; // @[LoadQueue.scala 163:19:@16229.4]
  wire  _T_16823; // @[LoadQueue.scala 163:13:@16230.4]
  wire  storeAddrNotKnownFlags_0_8; // @[LoadQueue.scala 163:19:@16231.4]
  wire  _T_16826; // @[LoadQueue.scala 163:13:@16232.4]
  wire  storeAddrNotKnownFlags_0_9; // @[LoadQueue.scala 163:19:@16233.4]
  wire  _T_16829; // @[LoadQueue.scala 163:13:@16234.4]
  wire  storeAddrNotKnownFlags_0_10; // @[LoadQueue.scala 163:19:@16235.4]
  wire  _T_16832; // @[LoadQueue.scala 163:13:@16236.4]
  wire  storeAddrNotKnownFlags_0_11; // @[LoadQueue.scala 163:19:@16237.4]
  wire  _T_16835; // @[LoadQueue.scala 163:13:@16238.4]
  wire  storeAddrNotKnownFlags_0_12; // @[LoadQueue.scala 163:19:@16239.4]
  wire  _T_16838; // @[LoadQueue.scala 163:13:@16240.4]
  wire  storeAddrNotKnownFlags_0_13; // @[LoadQueue.scala 163:19:@16241.4]
  wire  _T_16841; // @[LoadQueue.scala 163:13:@16242.4]
  wire  storeAddrNotKnownFlags_0_14; // @[LoadQueue.scala 163:19:@16243.4]
  wire  _T_16844; // @[LoadQueue.scala 163:13:@16244.4]
  wire  storeAddrNotKnownFlags_0_15; // @[LoadQueue.scala 163:19:@16245.4]
  wire  storeAddrNotKnownFlags_1_0; // @[LoadQueue.scala 163:19:@16263.4]
  wire  storeAddrNotKnownFlags_1_1; // @[LoadQueue.scala 163:19:@16265.4]
  wire  storeAddrNotKnownFlags_1_2; // @[LoadQueue.scala 163:19:@16267.4]
  wire  storeAddrNotKnownFlags_1_3; // @[LoadQueue.scala 163:19:@16269.4]
  wire  storeAddrNotKnownFlags_1_4; // @[LoadQueue.scala 163:19:@16271.4]
  wire  storeAddrNotKnownFlags_1_5; // @[LoadQueue.scala 163:19:@16273.4]
  wire  storeAddrNotKnownFlags_1_6; // @[LoadQueue.scala 163:19:@16275.4]
  wire  storeAddrNotKnownFlags_1_7; // @[LoadQueue.scala 163:19:@16277.4]
  wire  storeAddrNotKnownFlags_1_8; // @[LoadQueue.scala 163:19:@16279.4]
  wire  storeAddrNotKnownFlags_1_9; // @[LoadQueue.scala 163:19:@16281.4]
  wire  storeAddrNotKnownFlags_1_10; // @[LoadQueue.scala 163:19:@16283.4]
  wire  storeAddrNotKnownFlags_1_11; // @[LoadQueue.scala 163:19:@16285.4]
  wire  storeAddrNotKnownFlags_1_12; // @[LoadQueue.scala 163:19:@16287.4]
  wire  storeAddrNotKnownFlags_1_13; // @[LoadQueue.scala 163:19:@16289.4]
  wire  storeAddrNotKnownFlags_1_14; // @[LoadQueue.scala 163:19:@16291.4]
  wire  storeAddrNotKnownFlags_1_15; // @[LoadQueue.scala 163:19:@16293.4]
  wire  storeAddrNotKnownFlags_2_0; // @[LoadQueue.scala 163:19:@16311.4]
  wire  storeAddrNotKnownFlags_2_1; // @[LoadQueue.scala 163:19:@16313.4]
  wire  storeAddrNotKnownFlags_2_2; // @[LoadQueue.scala 163:19:@16315.4]
  wire  storeAddrNotKnownFlags_2_3; // @[LoadQueue.scala 163:19:@16317.4]
  wire  storeAddrNotKnownFlags_2_4; // @[LoadQueue.scala 163:19:@16319.4]
  wire  storeAddrNotKnownFlags_2_5; // @[LoadQueue.scala 163:19:@16321.4]
  wire  storeAddrNotKnownFlags_2_6; // @[LoadQueue.scala 163:19:@16323.4]
  wire  storeAddrNotKnownFlags_2_7; // @[LoadQueue.scala 163:19:@16325.4]
  wire  storeAddrNotKnownFlags_2_8; // @[LoadQueue.scala 163:19:@16327.4]
  wire  storeAddrNotKnownFlags_2_9; // @[LoadQueue.scala 163:19:@16329.4]
  wire  storeAddrNotKnownFlags_2_10; // @[LoadQueue.scala 163:19:@16331.4]
  wire  storeAddrNotKnownFlags_2_11; // @[LoadQueue.scala 163:19:@16333.4]
  wire  storeAddrNotKnownFlags_2_12; // @[LoadQueue.scala 163:19:@16335.4]
  wire  storeAddrNotKnownFlags_2_13; // @[LoadQueue.scala 163:19:@16337.4]
  wire  storeAddrNotKnownFlags_2_14; // @[LoadQueue.scala 163:19:@16339.4]
  wire  storeAddrNotKnownFlags_2_15; // @[LoadQueue.scala 163:19:@16341.4]
  wire  storeAddrNotKnownFlags_3_0; // @[LoadQueue.scala 163:19:@16359.4]
  wire  storeAddrNotKnownFlags_3_1; // @[LoadQueue.scala 163:19:@16361.4]
  wire  storeAddrNotKnownFlags_3_2; // @[LoadQueue.scala 163:19:@16363.4]
  wire  storeAddrNotKnownFlags_3_3; // @[LoadQueue.scala 163:19:@16365.4]
  wire  storeAddrNotKnownFlags_3_4; // @[LoadQueue.scala 163:19:@16367.4]
  wire  storeAddrNotKnownFlags_3_5; // @[LoadQueue.scala 163:19:@16369.4]
  wire  storeAddrNotKnownFlags_3_6; // @[LoadQueue.scala 163:19:@16371.4]
  wire  storeAddrNotKnownFlags_3_7; // @[LoadQueue.scala 163:19:@16373.4]
  wire  storeAddrNotKnownFlags_3_8; // @[LoadQueue.scala 163:19:@16375.4]
  wire  storeAddrNotKnownFlags_3_9; // @[LoadQueue.scala 163:19:@16377.4]
  wire  storeAddrNotKnownFlags_3_10; // @[LoadQueue.scala 163:19:@16379.4]
  wire  storeAddrNotKnownFlags_3_11; // @[LoadQueue.scala 163:19:@16381.4]
  wire  storeAddrNotKnownFlags_3_12; // @[LoadQueue.scala 163:19:@16383.4]
  wire  storeAddrNotKnownFlags_3_13; // @[LoadQueue.scala 163:19:@16385.4]
  wire  storeAddrNotKnownFlags_3_14; // @[LoadQueue.scala 163:19:@16387.4]
  wire  storeAddrNotKnownFlags_3_15; // @[LoadQueue.scala 163:19:@16389.4]
  wire  storeAddrNotKnownFlags_4_0; // @[LoadQueue.scala 163:19:@16407.4]
  wire  storeAddrNotKnownFlags_4_1; // @[LoadQueue.scala 163:19:@16409.4]
  wire  storeAddrNotKnownFlags_4_2; // @[LoadQueue.scala 163:19:@16411.4]
  wire  storeAddrNotKnownFlags_4_3; // @[LoadQueue.scala 163:19:@16413.4]
  wire  storeAddrNotKnownFlags_4_4; // @[LoadQueue.scala 163:19:@16415.4]
  wire  storeAddrNotKnownFlags_4_5; // @[LoadQueue.scala 163:19:@16417.4]
  wire  storeAddrNotKnownFlags_4_6; // @[LoadQueue.scala 163:19:@16419.4]
  wire  storeAddrNotKnownFlags_4_7; // @[LoadQueue.scala 163:19:@16421.4]
  wire  storeAddrNotKnownFlags_4_8; // @[LoadQueue.scala 163:19:@16423.4]
  wire  storeAddrNotKnownFlags_4_9; // @[LoadQueue.scala 163:19:@16425.4]
  wire  storeAddrNotKnownFlags_4_10; // @[LoadQueue.scala 163:19:@16427.4]
  wire  storeAddrNotKnownFlags_4_11; // @[LoadQueue.scala 163:19:@16429.4]
  wire  storeAddrNotKnownFlags_4_12; // @[LoadQueue.scala 163:19:@16431.4]
  wire  storeAddrNotKnownFlags_4_13; // @[LoadQueue.scala 163:19:@16433.4]
  wire  storeAddrNotKnownFlags_4_14; // @[LoadQueue.scala 163:19:@16435.4]
  wire  storeAddrNotKnownFlags_4_15; // @[LoadQueue.scala 163:19:@16437.4]
  wire  storeAddrNotKnownFlags_5_0; // @[LoadQueue.scala 163:19:@16455.4]
  wire  storeAddrNotKnownFlags_5_1; // @[LoadQueue.scala 163:19:@16457.4]
  wire  storeAddrNotKnownFlags_5_2; // @[LoadQueue.scala 163:19:@16459.4]
  wire  storeAddrNotKnownFlags_5_3; // @[LoadQueue.scala 163:19:@16461.4]
  wire  storeAddrNotKnownFlags_5_4; // @[LoadQueue.scala 163:19:@16463.4]
  wire  storeAddrNotKnownFlags_5_5; // @[LoadQueue.scala 163:19:@16465.4]
  wire  storeAddrNotKnownFlags_5_6; // @[LoadQueue.scala 163:19:@16467.4]
  wire  storeAddrNotKnownFlags_5_7; // @[LoadQueue.scala 163:19:@16469.4]
  wire  storeAddrNotKnownFlags_5_8; // @[LoadQueue.scala 163:19:@16471.4]
  wire  storeAddrNotKnownFlags_5_9; // @[LoadQueue.scala 163:19:@16473.4]
  wire  storeAddrNotKnownFlags_5_10; // @[LoadQueue.scala 163:19:@16475.4]
  wire  storeAddrNotKnownFlags_5_11; // @[LoadQueue.scala 163:19:@16477.4]
  wire  storeAddrNotKnownFlags_5_12; // @[LoadQueue.scala 163:19:@16479.4]
  wire  storeAddrNotKnownFlags_5_13; // @[LoadQueue.scala 163:19:@16481.4]
  wire  storeAddrNotKnownFlags_5_14; // @[LoadQueue.scala 163:19:@16483.4]
  wire  storeAddrNotKnownFlags_5_15; // @[LoadQueue.scala 163:19:@16485.4]
  wire  storeAddrNotKnownFlags_6_0; // @[LoadQueue.scala 163:19:@16503.4]
  wire  storeAddrNotKnownFlags_6_1; // @[LoadQueue.scala 163:19:@16505.4]
  wire  storeAddrNotKnownFlags_6_2; // @[LoadQueue.scala 163:19:@16507.4]
  wire  storeAddrNotKnownFlags_6_3; // @[LoadQueue.scala 163:19:@16509.4]
  wire  storeAddrNotKnownFlags_6_4; // @[LoadQueue.scala 163:19:@16511.4]
  wire  storeAddrNotKnownFlags_6_5; // @[LoadQueue.scala 163:19:@16513.4]
  wire  storeAddrNotKnownFlags_6_6; // @[LoadQueue.scala 163:19:@16515.4]
  wire  storeAddrNotKnownFlags_6_7; // @[LoadQueue.scala 163:19:@16517.4]
  wire  storeAddrNotKnownFlags_6_8; // @[LoadQueue.scala 163:19:@16519.4]
  wire  storeAddrNotKnownFlags_6_9; // @[LoadQueue.scala 163:19:@16521.4]
  wire  storeAddrNotKnownFlags_6_10; // @[LoadQueue.scala 163:19:@16523.4]
  wire  storeAddrNotKnownFlags_6_11; // @[LoadQueue.scala 163:19:@16525.4]
  wire  storeAddrNotKnownFlags_6_12; // @[LoadQueue.scala 163:19:@16527.4]
  wire  storeAddrNotKnownFlags_6_13; // @[LoadQueue.scala 163:19:@16529.4]
  wire  storeAddrNotKnownFlags_6_14; // @[LoadQueue.scala 163:19:@16531.4]
  wire  storeAddrNotKnownFlags_6_15; // @[LoadQueue.scala 163:19:@16533.4]
  wire  storeAddrNotKnownFlags_7_0; // @[LoadQueue.scala 163:19:@16551.4]
  wire  storeAddrNotKnownFlags_7_1; // @[LoadQueue.scala 163:19:@16553.4]
  wire  storeAddrNotKnownFlags_7_2; // @[LoadQueue.scala 163:19:@16555.4]
  wire  storeAddrNotKnownFlags_7_3; // @[LoadQueue.scala 163:19:@16557.4]
  wire  storeAddrNotKnownFlags_7_4; // @[LoadQueue.scala 163:19:@16559.4]
  wire  storeAddrNotKnownFlags_7_5; // @[LoadQueue.scala 163:19:@16561.4]
  wire  storeAddrNotKnownFlags_7_6; // @[LoadQueue.scala 163:19:@16563.4]
  wire  storeAddrNotKnownFlags_7_7; // @[LoadQueue.scala 163:19:@16565.4]
  wire  storeAddrNotKnownFlags_7_8; // @[LoadQueue.scala 163:19:@16567.4]
  wire  storeAddrNotKnownFlags_7_9; // @[LoadQueue.scala 163:19:@16569.4]
  wire  storeAddrNotKnownFlags_7_10; // @[LoadQueue.scala 163:19:@16571.4]
  wire  storeAddrNotKnownFlags_7_11; // @[LoadQueue.scala 163:19:@16573.4]
  wire  storeAddrNotKnownFlags_7_12; // @[LoadQueue.scala 163:19:@16575.4]
  wire  storeAddrNotKnownFlags_7_13; // @[LoadQueue.scala 163:19:@16577.4]
  wire  storeAddrNotKnownFlags_7_14; // @[LoadQueue.scala 163:19:@16579.4]
  wire  storeAddrNotKnownFlags_7_15; // @[LoadQueue.scala 163:19:@16581.4]
  wire  storeAddrNotKnownFlags_8_0; // @[LoadQueue.scala 163:19:@16599.4]
  wire  storeAddrNotKnownFlags_8_1; // @[LoadQueue.scala 163:19:@16601.4]
  wire  storeAddrNotKnownFlags_8_2; // @[LoadQueue.scala 163:19:@16603.4]
  wire  storeAddrNotKnownFlags_8_3; // @[LoadQueue.scala 163:19:@16605.4]
  wire  storeAddrNotKnownFlags_8_4; // @[LoadQueue.scala 163:19:@16607.4]
  wire  storeAddrNotKnownFlags_8_5; // @[LoadQueue.scala 163:19:@16609.4]
  wire  storeAddrNotKnownFlags_8_6; // @[LoadQueue.scala 163:19:@16611.4]
  wire  storeAddrNotKnownFlags_8_7; // @[LoadQueue.scala 163:19:@16613.4]
  wire  storeAddrNotKnownFlags_8_8; // @[LoadQueue.scala 163:19:@16615.4]
  wire  storeAddrNotKnownFlags_8_9; // @[LoadQueue.scala 163:19:@16617.4]
  wire  storeAddrNotKnownFlags_8_10; // @[LoadQueue.scala 163:19:@16619.4]
  wire  storeAddrNotKnownFlags_8_11; // @[LoadQueue.scala 163:19:@16621.4]
  wire  storeAddrNotKnownFlags_8_12; // @[LoadQueue.scala 163:19:@16623.4]
  wire  storeAddrNotKnownFlags_8_13; // @[LoadQueue.scala 163:19:@16625.4]
  wire  storeAddrNotKnownFlags_8_14; // @[LoadQueue.scala 163:19:@16627.4]
  wire  storeAddrNotKnownFlags_8_15; // @[LoadQueue.scala 163:19:@16629.4]
  wire  storeAddrNotKnownFlags_9_0; // @[LoadQueue.scala 163:19:@16647.4]
  wire  storeAddrNotKnownFlags_9_1; // @[LoadQueue.scala 163:19:@16649.4]
  wire  storeAddrNotKnownFlags_9_2; // @[LoadQueue.scala 163:19:@16651.4]
  wire  storeAddrNotKnownFlags_9_3; // @[LoadQueue.scala 163:19:@16653.4]
  wire  storeAddrNotKnownFlags_9_4; // @[LoadQueue.scala 163:19:@16655.4]
  wire  storeAddrNotKnownFlags_9_5; // @[LoadQueue.scala 163:19:@16657.4]
  wire  storeAddrNotKnownFlags_9_6; // @[LoadQueue.scala 163:19:@16659.4]
  wire  storeAddrNotKnownFlags_9_7; // @[LoadQueue.scala 163:19:@16661.4]
  wire  storeAddrNotKnownFlags_9_8; // @[LoadQueue.scala 163:19:@16663.4]
  wire  storeAddrNotKnownFlags_9_9; // @[LoadQueue.scala 163:19:@16665.4]
  wire  storeAddrNotKnownFlags_9_10; // @[LoadQueue.scala 163:19:@16667.4]
  wire  storeAddrNotKnownFlags_9_11; // @[LoadQueue.scala 163:19:@16669.4]
  wire  storeAddrNotKnownFlags_9_12; // @[LoadQueue.scala 163:19:@16671.4]
  wire  storeAddrNotKnownFlags_9_13; // @[LoadQueue.scala 163:19:@16673.4]
  wire  storeAddrNotKnownFlags_9_14; // @[LoadQueue.scala 163:19:@16675.4]
  wire  storeAddrNotKnownFlags_9_15; // @[LoadQueue.scala 163:19:@16677.4]
  wire  storeAddrNotKnownFlags_10_0; // @[LoadQueue.scala 163:19:@16695.4]
  wire  storeAddrNotKnownFlags_10_1; // @[LoadQueue.scala 163:19:@16697.4]
  wire  storeAddrNotKnownFlags_10_2; // @[LoadQueue.scala 163:19:@16699.4]
  wire  storeAddrNotKnownFlags_10_3; // @[LoadQueue.scala 163:19:@16701.4]
  wire  storeAddrNotKnownFlags_10_4; // @[LoadQueue.scala 163:19:@16703.4]
  wire  storeAddrNotKnownFlags_10_5; // @[LoadQueue.scala 163:19:@16705.4]
  wire  storeAddrNotKnownFlags_10_6; // @[LoadQueue.scala 163:19:@16707.4]
  wire  storeAddrNotKnownFlags_10_7; // @[LoadQueue.scala 163:19:@16709.4]
  wire  storeAddrNotKnownFlags_10_8; // @[LoadQueue.scala 163:19:@16711.4]
  wire  storeAddrNotKnownFlags_10_9; // @[LoadQueue.scala 163:19:@16713.4]
  wire  storeAddrNotKnownFlags_10_10; // @[LoadQueue.scala 163:19:@16715.4]
  wire  storeAddrNotKnownFlags_10_11; // @[LoadQueue.scala 163:19:@16717.4]
  wire  storeAddrNotKnownFlags_10_12; // @[LoadQueue.scala 163:19:@16719.4]
  wire  storeAddrNotKnownFlags_10_13; // @[LoadQueue.scala 163:19:@16721.4]
  wire  storeAddrNotKnownFlags_10_14; // @[LoadQueue.scala 163:19:@16723.4]
  wire  storeAddrNotKnownFlags_10_15; // @[LoadQueue.scala 163:19:@16725.4]
  wire  storeAddrNotKnownFlags_11_0; // @[LoadQueue.scala 163:19:@16743.4]
  wire  storeAddrNotKnownFlags_11_1; // @[LoadQueue.scala 163:19:@16745.4]
  wire  storeAddrNotKnownFlags_11_2; // @[LoadQueue.scala 163:19:@16747.4]
  wire  storeAddrNotKnownFlags_11_3; // @[LoadQueue.scala 163:19:@16749.4]
  wire  storeAddrNotKnownFlags_11_4; // @[LoadQueue.scala 163:19:@16751.4]
  wire  storeAddrNotKnownFlags_11_5; // @[LoadQueue.scala 163:19:@16753.4]
  wire  storeAddrNotKnownFlags_11_6; // @[LoadQueue.scala 163:19:@16755.4]
  wire  storeAddrNotKnownFlags_11_7; // @[LoadQueue.scala 163:19:@16757.4]
  wire  storeAddrNotKnownFlags_11_8; // @[LoadQueue.scala 163:19:@16759.4]
  wire  storeAddrNotKnownFlags_11_9; // @[LoadQueue.scala 163:19:@16761.4]
  wire  storeAddrNotKnownFlags_11_10; // @[LoadQueue.scala 163:19:@16763.4]
  wire  storeAddrNotKnownFlags_11_11; // @[LoadQueue.scala 163:19:@16765.4]
  wire  storeAddrNotKnownFlags_11_12; // @[LoadQueue.scala 163:19:@16767.4]
  wire  storeAddrNotKnownFlags_11_13; // @[LoadQueue.scala 163:19:@16769.4]
  wire  storeAddrNotKnownFlags_11_14; // @[LoadQueue.scala 163:19:@16771.4]
  wire  storeAddrNotKnownFlags_11_15; // @[LoadQueue.scala 163:19:@16773.4]
  wire  storeAddrNotKnownFlags_12_0; // @[LoadQueue.scala 163:19:@16791.4]
  wire  storeAddrNotKnownFlags_12_1; // @[LoadQueue.scala 163:19:@16793.4]
  wire  storeAddrNotKnownFlags_12_2; // @[LoadQueue.scala 163:19:@16795.4]
  wire  storeAddrNotKnownFlags_12_3; // @[LoadQueue.scala 163:19:@16797.4]
  wire  storeAddrNotKnownFlags_12_4; // @[LoadQueue.scala 163:19:@16799.4]
  wire  storeAddrNotKnownFlags_12_5; // @[LoadQueue.scala 163:19:@16801.4]
  wire  storeAddrNotKnownFlags_12_6; // @[LoadQueue.scala 163:19:@16803.4]
  wire  storeAddrNotKnownFlags_12_7; // @[LoadQueue.scala 163:19:@16805.4]
  wire  storeAddrNotKnownFlags_12_8; // @[LoadQueue.scala 163:19:@16807.4]
  wire  storeAddrNotKnownFlags_12_9; // @[LoadQueue.scala 163:19:@16809.4]
  wire  storeAddrNotKnownFlags_12_10; // @[LoadQueue.scala 163:19:@16811.4]
  wire  storeAddrNotKnownFlags_12_11; // @[LoadQueue.scala 163:19:@16813.4]
  wire  storeAddrNotKnownFlags_12_12; // @[LoadQueue.scala 163:19:@16815.4]
  wire  storeAddrNotKnownFlags_12_13; // @[LoadQueue.scala 163:19:@16817.4]
  wire  storeAddrNotKnownFlags_12_14; // @[LoadQueue.scala 163:19:@16819.4]
  wire  storeAddrNotKnownFlags_12_15; // @[LoadQueue.scala 163:19:@16821.4]
  wire  storeAddrNotKnownFlags_13_0; // @[LoadQueue.scala 163:19:@16839.4]
  wire  storeAddrNotKnownFlags_13_1; // @[LoadQueue.scala 163:19:@16841.4]
  wire  storeAddrNotKnownFlags_13_2; // @[LoadQueue.scala 163:19:@16843.4]
  wire  storeAddrNotKnownFlags_13_3; // @[LoadQueue.scala 163:19:@16845.4]
  wire  storeAddrNotKnownFlags_13_4; // @[LoadQueue.scala 163:19:@16847.4]
  wire  storeAddrNotKnownFlags_13_5; // @[LoadQueue.scala 163:19:@16849.4]
  wire  storeAddrNotKnownFlags_13_6; // @[LoadQueue.scala 163:19:@16851.4]
  wire  storeAddrNotKnownFlags_13_7; // @[LoadQueue.scala 163:19:@16853.4]
  wire  storeAddrNotKnownFlags_13_8; // @[LoadQueue.scala 163:19:@16855.4]
  wire  storeAddrNotKnownFlags_13_9; // @[LoadQueue.scala 163:19:@16857.4]
  wire  storeAddrNotKnownFlags_13_10; // @[LoadQueue.scala 163:19:@16859.4]
  wire  storeAddrNotKnownFlags_13_11; // @[LoadQueue.scala 163:19:@16861.4]
  wire  storeAddrNotKnownFlags_13_12; // @[LoadQueue.scala 163:19:@16863.4]
  wire  storeAddrNotKnownFlags_13_13; // @[LoadQueue.scala 163:19:@16865.4]
  wire  storeAddrNotKnownFlags_13_14; // @[LoadQueue.scala 163:19:@16867.4]
  wire  storeAddrNotKnownFlags_13_15; // @[LoadQueue.scala 163:19:@16869.4]
  wire  storeAddrNotKnownFlags_14_0; // @[LoadQueue.scala 163:19:@16887.4]
  wire  storeAddrNotKnownFlags_14_1; // @[LoadQueue.scala 163:19:@16889.4]
  wire  storeAddrNotKnownFlags_14_2; // @[LoadQueue.scala 163:19:@16891.4]
  wire  storeAddrNotKnownFlags_14_3; // @[LoadQueue.scala 163:19:@16893.4]
  wire  storeAddrNotKnownFlags_14_4; // @[LoadQueue.scala 163:19:@16895.4]
  wire  storeAddrNotKnownFlags_14_5; // @[LoadQueue.scala 163:19:@16897.4]
  wire  storeAddrNotKnownFlags_14_6; // @[LoadQueue.scala 163:19:@16899.4]
  wire  storeAddrNotKnownFlags_14_7; // @[LoadQueue.scala 163:19:@16901.4]
  wire  storeAddrNotKnownFlags_14_8; // @[LoadQueue.scala 163:19:@16903.4]
  wire  storeAddrNotKnownFlags_14_9; // @[LoadQueue.scala 163:19:@16905.4]
  wire  storeAddrNotKnownFlags_14_10; // @[LoadQueue.scala 163:19:@16907.4]
  wire  storeAddrNotKnownFlags_14_11; // @[LoadQueue.scala 163:19:@16909.4]
  wire  storeAddrNotKnownFlags_14_12; // @[LoadQueue.scala 163:19:@16911.4]
  wire  storeAddrNotKnownFlags_14_13; // @[LoadQueue.scala 163:19:@16913.4]
  wire  storeAddrNotKnownFlags_14_14; // @[LoadQueue.scala 163:19:@16915.4]
  wire  storeAddrNotKnownFlags_14_15; // @[LoadQueue.scala 163:19:@16917.4]
  wire  storeAddrNotKnownFlags_15_0; // @[LoadQueue.scala 163:19:@16935.4]
  wire  storeAddrNotKnownFlags_15_1; // @[LoadQueue.scala 163:19:@16937.4]
  wire  storeAddrNotKnownFlags_15_2; // @[LoadQueue.scala 163:19:@16939.4]
  wire  storeAddrNotKnownFlags_15_3; // @[LoadQueue.scala 163:19:@16941.4]
  wire  storeAddrNotKnownFlags_15_4; // @[LoadQueue.scala 163:19:@16943.4]
  wire  storeAddrNotKnownFlags_15_5; // @[LoadQueue.scala 163:19:@16945.4]
  wire  storeAddrNotKnownFlags_15_6; // @[LoadQueue.scala 163:19:@16947.4]
  wire  storeAddrNotKnownFlags_15_7; // @[LoadQueue.scala 163:19:@16949.4]
  wire  storeAddrNotKnownFlags_15_8; // @[LoadQueue.scala 163:19:@16951.4]
  wire  storeAddrNotKnownFlags_15_9; // @[LoadQueue.scala 163:19:@16953.4]
  wire  storeAddrNotKnownFlags_15_10; // @[LoadQueue.scala 163:19:@16955.4]
  wire  storeAddrNotKnownFlags_15_11; // @[LoadQueue.scala 163:19:@16957.4]
  wire  storeAddrNotKnownFlags_15_12; // @[LoadQueue.scala 163:19:@16959.4]
  wire  storeAddrNotKnownFlags_15_13; // @[LoadQueue.scala 163:19:@16961.4]
  wire  storeAddrNotKnownFlags_15_14; // @[LoadQueue.scala 163:19:@16963.4]
  wire  storeAddrNotKnownFlags_15_15; // @[LoadQueue.scala 163:19:@16965.4]
  wire [7:0] _T_18002; // @[Mux.scala 19:72:@17296.4]
  wire [7:0] _T_18009; // @[Mux.scala 19:72:@17303.4]
  wire [15:0] _T_18010; // @[Mux.scala 19:72:@17304.4]
  wire [15:0] _T_18012; // @[Mux.scala 19:72:@17305.4]
  wire [7:0] _T_18019; // @[Mux.scala 19:72:@17312.4]
  wire [7:0] _T_18026; // @[Mux.scala 19:72:@17319.4]
  wire [15:0] _T_18027; // @[Mux.scala 19:72:@17320.4]
  wire [15:0] _T_18029; // @[Mux.scala 19:72:@17321.4]
  wire [7:0] _T_18036; // @[Mux.scala 19:72:@17328.4]
  wire [7:0] _T_18043; // @[Mux.scala 19:72:@17335.4]
  wire [15:0] _T_18044; // @[Mux.scala 19:72:@17336.4]
  wire [15:0] _T_18046; // @[Mux.scala 19:72:@17337.4]
  wire [7:0] _T_18053; // @[Mux.scala 19:72:@17344.4]
  wire [7:0] _T_18060; // @[Mux.scala 19:72:@17351.4]
  wire [15:0] _T_18061; // @[Mux.scala 19:72:@17352.4]
  wire [15:0] _T_18063; // @[Mux.scala 19:72:@17353.4]
  wire [7:0] _T_18070; // @[Mux.scala 19:72:@17360.4]
  wire [7:0] _T_18077; // @[Mux.scala 19:72:@17367.4]
  wire [15:0] _T_18078; // @[Mux.scala 19:72:@17368.4]
  wire [15:0] _T_18080; // @[Mux.scala 19:72:@17369.4]
  wire [7:0] _T_18087; // @[Mux.scala 19:72:@17376.4]
  wire [7:0] _T_18094; // @[Mux.scala 19:72:@17383.4]
  wire [15:0] _T_18095; // @[Mux.scala 19:72:@17384.4]
  wire [15:0] _T_18097; // @[Mux.scala 19:72:@17385.4]
  wire [7:0] _T_18104; // @[Mux.scala 19:72:@17392.4]
  wire [7:0] _T_18111; // @[Mux.scala 19:72:@17399.4]
  wire [15:0] _T_18112; // @[Mux.scala 19:72:@17400.4]
  wire [15:0] _T_18114; // @[Mux.scala 19:72:@17401.4]
  wire [7:0] _T_18121; // @[Mux.scala 19:72:@17408.4]
  wire [7:0] _T_18128; // @[Mux.scala 19:72:@17415.4]
  wire [15:0] _T_18129; // @[Mux.scala 19:72:@17416.4]
  wire [15:0] _T_18131; // @[Mux.scala 19:72:@17417.4]
  wire [15:0] _T_18146; // @[Mux.scala 19:72:@17432.4]
  wire [15:0] _T_18148; // @[Mux.scala 19:72:@17433.4]
  wire [15:0] _T_18163; // @[Mux.scala 19:72:@17448.4]
  wire [15:0] _T_18165; // @[Mux.scala 19:72:@17449.4]
  wire [15:0] _T_18180; // @[Mux.scala 19:72:@17464.4]
  wire [15:0] _T_18182; // @[Mux.scala 19:72:@17465.4]
  wire [15:0] _T_18197; // @[Mux.scala 19:72:@17480.4]
  wire [15:0] _T_18199; // @[Mux.scala 19:72:@17481.4]
  wire [15:0] _T_18214; // @[Mux.scala 19:72:@17496.4]
  wire [15:0] _T_18216; // @[Mux.scala 19:72:@17497.4]
  wire [15:0] _T_18231; // @[Mux.scala 19:72:@17512.4]
  wire [15:0] _T_18233; // @[Mux.scala 19:72:@17513.4]
  wire [15:0] _T_18248; // @[Mux.scala 19:72:@17528.4]
  wire [15:0] _T_18250; // @[Mux.scala 19:72:@17529.4]
  wire [15:0] _T_18265; // @[Mux.scala 19:72:@17544.4]
  wire [15:0] _T_18267; // @[Mux.scala 19:72:@17545.4]
  wire [15:0] _T_18268; // @[Mux.scala 19:72:@17546.4]
  wire [15:0] _T_18269; // @[Mux.scala 19:72:@17547.4]
  wire [15:0] _T_18270; // @[Mux.scala 19:72:@17548.4]
  wire [15:0] _T_18271; // @[Mux.scala 19:72:@17549.4]
  wire [15:0] _T_18272; // @[Mux.scala 19:72:@17550.4]
  wire [15:0] _T_18273; // @[Mux.scala 19:72:@17551.4]
  wire [15:0] _T_18274; // @[Mux.scala 19:72:@17552.4]
  wire [15:0] _T_18275; // @[Mux.scala 19:72:@17553.4]
  wire [15:0] _T_18276; // @[Mux.scala 19:72:@17554.4]
  wire [15:0] _T_18277; // @[Mux.scala 19:72:@17555.4]
  wire [15:0] _T_18278; // @[Mux.scala 19:72:@17556.4]
  wire [15:0] _T_18279; // @[Mux.scala 19:72:@17557.4]
  wire [15:0] _T_18280; // @[Mux.scala 19:72:@17558.4]
  wire [15:0] _T_18281; // @[Mux.scala 19:72:@17559.4]
  wire [15:0] _T_18282; // @[Mux.scala 19:72:@17560.4]
  wire [7:0] _T_18860; // @[Mux.scala 19:72:@17910.4]
  wire [7:0] _T_18867; // @[Mux.scala 19:72:@17917.4]
  wire [15:0] _T_18868; // @[Mux.scala 19:72:@17918.4]
  wire [15:0] _T_18870; // @[Mux.scala 19:72:@17919.4]
  wire [7:0] _T_18877; // @[Mux.scala 19:72:@17926.4]
  wire [7:0] _T_18884; // @[Mux.scala 19:72:@17933.4]
  wire [15:0] _T_18885; // @[Mux.scala 19:72:@17934.4]
  wire [15:0] _T_18887; // @[Mux.scala 19:72:@17935.4]
  wire [7:0] _T_18894; // @[Mux.scala 19:72:@17942.4]
  wire [7:0] _T_18901; // @[Mux.scala 19:72:@17949.4]
  wire [15:0] _T_18902; // @[Mux.scala 19:72:@17950.4]
  wire [15:0] _T_18904; // @[Mux.scala 19:72:@17951.4]
  wire [7:0] _T_18911; // @[Mux.scala 19:72:@17958.4]
  wire [7:0] _T_18918; // @[Mux.scala 19:72:@17965.4]
  wire [15:0] _T_18919; // @[Mux.scala 19:72:@17966.4]
  wire [15:0] _T_18921; // @[Mux.scala 19:72:@17967.4]
  wire [7:0] _T_18928; // @[Mux.scala 19:72:@17974.4]
  wire [7:0] _T_18935; // @[Mux.scala 19:72:@17981.4]
  wire [15:0] _T_18936; // @[Mux.scala 19:72:@17982.4]
  wire [15:0] _T_18938; // @[Mux.scala 19:72:@17983.4]
  wire [7:0] _T_18945; // @[Mux.scala 19:72:@17990.4]
  wire [7:0] _T_18952; // @[Mux.scala 19:72:@17997.4]
  wire [15:0] _T_18953; // @[Mux.scala 19:72:@17998.4]
  wire [15:0] _T_18955; // @[Mux.scala 19:72:@17999.4]
  wire [7:0] _T_18962; // @[Mux.scala 19:72:@18006.4]
  wire [7:0] _T_18969; // @[Mux.scala 19:72:@18013.4]
  wire [15:0] _T_18970; // @[Mux.scala 19:72:@18014.4]
  wire [15:0] _T_18972; // @[Mux.scala 19:72:@18015.4]
  wire [7:0] _T_18979; // @[Mux.scala 19:72:@18022.4]
  wire [7:0] _T_18986; // @[Mux.scala 19:72:@18029.4]
  wire [15:0] _T_18987; // @[Mux.scala 19:72:@18030.4]
  wire [15:0] _T_18989; // @[Mux.scala 19:72:@18031.4]
  wire [15:0] _T_19004; // @[Mux.scala 19:72:@18046.4]
  wire [15:0] _T_19006; // @[Mux.scala 19:72:@18047.4]
  wire [15:0] _T_19021; // @[Mux.scala 19:72:@18062.4]
  wire [15:0] _T_19023; // @[Mux.scala 19:72:@18063.4]
  wire [15:0] _T_19038; // @[Mux.scala 19:72:@18078.4]
  wire [15:0] _T_19040; // @[Mux.scala 19:72:@18079.4]
  wire [15:0] _T_19055; // @[Mux.scala 19:72:@18094.4]
  wire [15:0] _T_19057; // @[Mux.scala 19:72:@18095.4]
  wire [15:0] _T_19072; // @[Mux.scala 19:72:@18110.4]
  wire [15:0] _T_19074; // @[Mux.scala 19:72:@18111.4]
  wire [15:0] _T_19089; // @[Mux.scala 19:72:@18126.4]
  wire [15:0] _T_19091; // @[Mux.scala 19:72:@18127.4]
  wire [15:0] _T_19106; // @[Mux.scala 19:72:@18142.4]
  wire [15:0] _T_19108; // @[Mux.scala 19:72:@18143.4]
  wire [15:0] _T_19123; // @[Mux.scala 19:72:@18158.4]
  wire [15:0] _T_19125; // @[Mux.scala 19:72:@18159.4]
  wire [15:0] _T_19126; // @[Mux.scala 19:72:@18160.4]
  wire [15:0] _T_19127; // @[Mux.scala 19:72:@18161.4]
  wire [15:0] _T_19128; // @[Mux.scala 19:72:@18162.4]
  wire [15:0] _T_19129; // @[Mux.scala 19:72:@18163.4]
  wire [15:0] _T_19130; // @[Mux.scala 19:72:@18164.4]
  wire [15:0] _T_19131; // @[Mux.scala 19:72:@18165.4]
  wire [15:0] _T_19132; // @[Mux.scala 19:72:@18166.4]
  wire [15:0] _T_19133; // @[Mux.scala 19:72:@18167.4]
  wire [15:0] _T_19134; // @[Mux.scala 19:72:@18168.4]
  wire [15:0] _T_19135; // @[Mux.scala 19:72:@18169.4]
  wire [15:0] _T_19136; // @[Mux.scala 19:72:@18170.4]
  wire [15:0] _T_19137; // @[Mux.scala 19:72:@18171.4]
  wire [15:0] _T_19138; // @[Mux.scala 19:72:@18172.4]
  wire [15:0] _T_19139; // @[Mux.scala 19:72:@18173.4]
  wire [15:0] _T_19140; // @[Mux.scala 19:72:@18174.4]
  wire [7:0] _T_19718; // @[Mux.scala 19:72:@18524.4]
  wire [7:0] _T_19725; // @[Mux.scala 19:72:@18531.4]
  wire [15:0] _T_19726; // @[Mux.scala 19:72:@18532.4]
  wire [15:0] _T_19728; // @[Mux.scala 19:72:@18533.4]
  wire [7:0] _T_19735; // @[Mux.scala 19:72:@18540.4]
  wire [7:0] _T_19742; // @[Mux.scala 19:72:@18547.4]
  wire [15:0] _T_19743; // @[Mux.scala 19:72:@18548.4]
  wire [15:0] _T_19745; // @[Mux.scala 19:72:@18549.4]
  wire [7:0] _T_19752; // @[Mux.scala 19:72:@18556.4]
  wire [7:0] _T_19759; // @[Mux.scala 19:72:@18563.4]
  wire [15:0] _T_19760; // @[Mux.scala 19:72:@18564.4]
  wire [15:0] _T_19762; // @[Mux.scala 19:72:@18565.4]
  wire [7:0] _T_19769; // @[Mux.scala 19:72:@18572.4]
  wire [7:0] _T_19776; // @[Mux.scala 19:72:@18579.4]
  wire [15:0] _T_19777; // @[Mux.scala 19:72:@18580.4]
  wire [15:0] _T_19779; // @[Mux.scala 19:72:@18581.4]
  wire [7:0] _T_19786; // @[Mux.scala 19:72:@18588.4]
  wire [7:0] _T_19793; // @[Mux.scala 19:72:@18595.4]
  wire [15:0] _T_19794; // @[Mux.scala 19:72:@18596.4]
  wire [15:0] _T_19796; // @[Mux.scala 19:72:@18597.4]
  wire [7:0] _T_19803; // @[Mux.scala 19:72:@18604.4]
  wire [7:0] _T_19810; // @[Mux.scala 19:72:@18611.4]
  wire [15:0] _T_19811; // @[Mux.scala 19:72:@18612.4]
  wire [15:0] _T_19813; // @[Mux.scala 19:72:@18613.4]
  wire [7:0] _T_19820; // @[Mux.scala 19:72:@18620.4]
  wire [7:0] _T_19827; // @[Mux.scala 19:72:@18627.4]
  wire [15:0] _T_19828; // @[Mux.scala 19:72:@18628.4]
  wire [15:0] _T_19830; // @[Mux.scala 19:72:@18629.4]
  wire [7:0] _T_19837; // @[Mux.scala 19:72:@18636.4]
  wire [7:0] _T_19844; // @[Mux.scala 19:72:@18643.4]
  wire [15:0] _T_19845; // @[Mux.scala 19:72:@18644.4]
  wire [15:0] _T_19847; // @[Mux.scala 19:72:@18645.4]
  wire [15:0] _T_19862; // @[Mux.scala 19:72:@18660.4]
  wire [15:0] _T_19864; // @[Mux.scala 19:72:@18661.4]
  wire [15:0] _T_19879; // @[Mux.scala 19:72:@18676.4]
  wire [15:0] _T_19881; // @[Mux.scala 19:72:@18677.4]
  wire [15:0] _T_19896; // @[Mux.scala 19:72:@18692.4]
  wire [15:0] _T_19898; // @[Mux.scala 19:72:@18693.4]
  wire [15:0] _T_19913; // @[Mux.scala 19:72:@18708.4]
  wire [15:0] _T_19915; // @[Mux.scala 19:72:@18709.4]
  wire [15:0] _T_19930; // @[Mux.scala 19:72:@18724.4]
  wire [15:0] _T_19932; // @[Mux.scala 19:72:@18725.4]
  wire [15:0] _T_19947; // @[Mux.scala 19:72:@18740.4]
  wire [15:0] _T_19949; // @[Mux.scala 19:72:@18741.4]
  wire [15:0] _T_19964; // @[Mux.scala 19:72:@18756.4]
  wire [15:0] _T_19966; // @[Mux.scala 19:72:@18757.4]
  wire [15:0] _T_19981; // @[Mux.scala 19:72:@18772.4]
  wire [15:0] _T_19983; // @[Mux.scala 19:72:@18773.4]
  wire [15:0] _T_19984; // @[Mux.scala 19:72:@18774.4]
  wire [15:0] _T_19985; // @[Mux.scala 19:72:@18775.4]
  wire [15:0] _T_19986; // @[Mux.scala 19:72:@18776.4]
  wire [15:0] _T_19987; // @[Mux.scala 19:72:@18777.4]
  wire [15:0] _T_19988; // @[Mux.scala 19:72:@18778.4]
  wire [15:0] _T_19989; // @[Mux.scala 19:72:@18779.4]
  wire [15:0] _T_19990; // @[Mux.scala 19:72:@18780.4]
  wire [15:0] _T_19991; // @[Mux.scala 19:72:@18781.4]
  wire [15:0] _T_19992; // @[Mux.scala 19:72:@18782.4]
  wire [15:0] _T_19993; // @[Mux.scala 19:72:@18783.4]
  wire [15:0] _T_19994; // @[Mux.scala 19:72:@18784.4]
  wire [15:0] _T_19995; // @[Mux.scala 19:72:@18785.4]
  wire [15:0] _T_19996; // @[Mux.scala 19:72:@18786.4]
  wire [15:0] _T_19997; // @[Mux.scala 19:72:@18787.4]
  wire [15:0] _T_19998; // @[Mux.scala 19:72:@18788.4]
  wire [7:0] _T_20576; // @[Mux.scala 19:72:@19138.4]
  wire [7:0] _T_20583; // @[Mux.scala 19:72:@19145.4]
  wire [15:0] _T_20584; // @[Mux.scala 19:72:@19146.4]
  wire [15:0] _T_20586; // @[Mux.scala 19:72:@19147.4]
  wire [7:0] _T_20593; // @[Mux.scala 19:72:@19154.4]
  wire [7:0] _T_20600; // @[Mux.scala 19:72:@19161.4]
  wire [15:0] _T_20601; // @[Mux.scala 19:72:@19162.4]
  wire [15:0] _T_20603; // @[Mux.scala 19:72:@19163.4]
  wire [7:0] _T_20610; // @[Mux.scala 19:72:@19170.4]
  wire [7:0] _T_20617; // @[Mux.scala 19:72:@19177.4]
  wire [15:0] _T_20618; // @[Mux.scala 19:72:@19178.4]
  wire [15:0] _T_20620; // @[Mux.scala 19:72:@19179.4]
  wire [7:0] _T_20627; // @[Mux.scala 19:72:@19186.4]
  wire [7:0] _T_20634; // @[Mux.scala 19:72:@19193.4]
  wire [15:0] _T_20635; // @[Mux.scala 19:72:@19194.4]
  wire [15:0] _T_20637; // @[Mux.scala 19:72:@19195.4]
  wire [7:0] _T_20644; // @[Mux.scala 19:72:@19202.4]
  wire [7:0] _T_20651; // @[Mux.scala 19:72:@19209.4]
  wire [15:0] _T_20652; // @[Mux.scala 19:72:@19210.4]
  wire [15:0] _T_20654; // @[Mux.scala 19:72:@19211.4]
  wire [7:0] _T_20661; // @[Mux.scala 19:72:@19218.4]
  wire [7:0] _T_20668; // @[Mux.scala 19:72:@19225.4]
  wire [15:0] _T_20669; // @[Mux.scala 19:72:@19226.4]
  wire [15:0] _T_20671; // @[Mux.scala 19:72:@19227.4]
  wire [7:0] _T_20678; // @[Mux.scala 19:72:@19234.4]
  wire [7:0] _T_20685; // @[Mux.scala 19:72:@19241.4]
  wire [15:0] _T_20686; // @[Mux.scala 19:72:@19242.4]
  wire [15:0] _T_20688; // @[Mux.scala 19:72:@19243.4]
  wire [7:0] _T_20695; // @[Mux.scala 19:72:@19250.4]
  wire [7:0] _T_20702; // @[Mux.scala 19:72:@19257.4]
  wire [15:0] _T_20703; // @[Mux.scala 19:72:@19258.4]
  wire [15:0] _T_20705; // @[Mux.scala 19:72:@19259.4]
  wire [15:0] _T_20720; // @[Mux.scala 19:72:@19274.4]
  wire [15:0] _T_20722; // @[Mux.scala 19:72:@19275.4]
  wire [15:0] _T_20737; // @[Mux.scala 19:72:@19290.4]
  wire [15:0] _T_20739; // @[Mux.scala 19:72:@19291.4]
  wire [15:0] _T_20754; // @[Mux.scala 19:72:@19306.4]
  wire [15:0] _T_20756; // @[Mux.scala 19:72:@19307.4]
  wire [15:0] _T_20771; // @[Mux.scala 19:72:@19322.4]
  wire [15:0] _T_20773; // @[Mux.scala 19:72:@19323.4]
  wire [15:0] _T_20788; // @[Mux.scala 19:72:@19338.4]
  wire [15:0] _T_20790; // @[Mux.scala 19:72:@19339.4]
  wire [15:0] _T_20805; // @[Mux.scala 19:72:@19354.4]
  wire [15:0] _T_20807; // @[Mux.scala 19:72:@19355.4]
  wire [15:0] _T_20822; // @[Mux.scala 19:72:@19370.4]
  wire [15:0] _T_20824; // @[Mux.scala 19:72:@19371.4]
  wire [15:0] _T_20839; // @[Mux.scala 19:72:@19386.4]
  wire [15:0] _T_20841; // @[Mux.scala 19:72:@19387.4]
  wire [15:0] _T_20842; // @[Mux.scala 19:72:@19388.4]
  wire [15:0] _T_20843; // @[Mux.scala 19:72:@19389.4]
  wire [15:0] _T_20844; // @[Mux.scala 19:72:@19390.4]
  wire [15:0] _T_20845; // @[Mux.scala 19:72:@19391.4]
  wire [15:0] _T_20846; // @[Mux.scala 19:72:@19392.4]
  wire [15:0] _T_20847; // @[Mux.scala 19:72:@19393.4]
  wire [15:0] _T_20848; // @[Mux.scala 19:72:@19394.4]
  wire [15:0] _T_20849; // @[Mux.scala 19:72:@19395.4]
  wire [15:0] _T_20850; // @[Mux.scala 19:72:@19396.4]
  wire [15:0] _T_20851; // @[Mux.scala 19:72:@19397.4]
  wire [15:0] _T_20852; // @[Mux.scala 19:72:@19398.4]
  wire [15:0] _T_20853; // @[Mux.scala 19:72:@19399.4]
  wire [15:0] _T_20854; // @[Mux.scala 19:72:@19400.4]
  wire [15:0] _T_20855; // @[Mux.scala 19:72:@19401.4]
  wire [15:0] _T_20856; // @[Mux.scala 19:72:@19402.4]
  wire [7:0] _T_21434; // @[Mux.scala 19:72:@19752.4]
  wire [7:0] _T_21441; // @[Mux.scala 19:72:@19759.4]
  wire [15:0] _T_21442; // @[Mux.scala 19:72:@19760.4]
  wire [15:0] _T_21444; // @[Mux.scala 19:72:@19761.4]
  wire [7:0] _T_21451; // @[Mux.scala 19:72:@19768.4]
  wire [7:0] _T_21458; // @[Mux.scala 19:72:@19775.4]
  wire [15:0] _T_21459; // @[Mux.scala 19:72:@19776.4]
  wire [15:0] _T_21461; // @[Mux.scala 19:72:@19777.4]
  wire [7:0] _T_21468; // @[Mux.scala 19:72:@19784.4]
  wire [7:0] _T_21475; // @[Mux.scala 19:72:@19791.4]
  wire [15:0] _T_21476; // @[Mux.scala 19:72:@19792.4]
  wire [15:0] _T_21478; // @[Mux.scala 19:72:@19793.4]
  wire [7:0] _T_21485; // @[Mux.scala 19:72:@19800.4]
  wire [7:0] _T_21492; // @[Mux.scala 19:72:@19807.4]
  wire [15:0] _T_21493; // @[Mux.scala 19:72:@19808.4]
  wire [15:0] _T_21495; // @[Mux.scala 19:72:@19809.4]
  wire [7:0] _T_21502; // @[Mux.scala 19:72:@19816.4]
  wire [7:0] _T_21509; // @[Mux.scala 19:72:@19823.4]
  wire [15:0] _T_21510; // @[Mux.scala 19:72:@19824.4]
  wire [15:0] _T_21512; // @[Mux.scala 19:72:@19825.4]
  wire [7:0] _T_21519; // @[Mux.scala 19:72:@19832.4]
  wire [7:0] _T_21526; // @[Mux.scala 19:72:@19839.4]
  wire [15:0] _T_21527; // @[Mux.scala 19:72:@19840.4]
  wire [15:0] _T_21529; // @[Mux.scala 19:72:@19841.4]
  wire [7:0] _T_21536; // @[Mux.scala 19:72:@19848.4]
  wire [7:0] _T_21543; // @[Mux.scala 19:72:@19855.4]
  wire [15:0] _T_21544; // @[Mux.scala 19:72:@19856.4]
  wire [15:0] _T_21546; // @[Mux.scala 19:72:@19857.4]
  wire [7:0] _T_21553; // @[Mux.scala 19:72:@19864.4]
  wire [7:0] _T_21560; // @[Mux.scala 19:72:@19871.4]
  wire [15:0] _T_21561; // @[Mux.scala 19:72:@19872.4]
  wire [15:0] _T_21563; // @[Mux.scala 19:72:@19873.4]
  wire [15:0] _T_21578; // @[Mux.scala 19:72:@19888.4]
  wire [15:0] _T_21580; // @[Mux.scala 19:72:@19889.4]
  wire [15:0] _T_21595; // @[Mux.scala 19:72:@19904.4]
  wire [15:0] _T_21597; // @[Mux.scala 19:72:@19905.4]
  wire [15:0] _T_21612; // @[Mux.scala 19:72:@19920.4]
  wire [15:0] _T_21614; // @[Mux.scala 19:72:@19921.4]
  wire [15:0] _T_21629; // @[Mux.scala 19:72:@19936.4]
  wire [15:0] _T_21631; // @[Mux.scala 19:72:@19937.4]
  wire [15:0] _T_21646; // @[Mux.scala 19:72:@19952.4]
  wire [15:0] _T_21648; // @[Mux.scala 19:72:@19953.4]
  wire [15:0] _T_21663; // @[Mux.scala 19:72:@19968.4]
  wire [15:0] _T_21665; // @[Mux.scala 19:72:@19969.4]
  wire [15:0] _T_21680; // @[Mux.scala 19:72:@19984.4]
  wire [15:0] _T_21682; // @[Mux.scala 19:72:@19985.4]
  wire [15:0] _T_21697; // @[Mux.scala 19:72:@20000.4]
  wire [15:0] _T_21699; // @[Mux.scala 19:72:@20001.4]
  wire [15:0] _T_21700; // @[Mux.scala 19:72:@20002.4]
  wire [15:0] _T_21701; // @[Mux.scala 19:72:@20003.4]
  wire [15:0] _T_21702; // @[Mux.scala 19:72:@20004.4]
  wire [15:0] _T_21703; // @[Mux.scala 19:72:@20005.4]
  wire [15:0] _T_21704; // @[Mux.scala 19:72:@20006.4]
  wire [15:0] _T_21705; // @[Mux.scala 19:72:@20007.4]
  wire [15:0] _T_21706; // @[Mux.scala 19:72:@20008.4]
  wire [15:0] _T_21707; // @[Mux.scala 19:72:@20009.4]
  wire [15:0] _T_21708; // @[Mux.scala 19:72:@20010.4]
  wire [15:0] _T_21709; // @[Mux.scala 19:72:@20011.4]
  wire [15:0] _T_21710; // @[Mux.scala 19:72:@20012.4]
  wire [15:0] _T_21711; // @[Mux.scala 19:72:@20013.4]
  wire [15:0] _T_21712; // @[Mux.scala 19:72:@20014.4]
  wire [15:0] _T_21713; // @[Mux.scala 19:72:@20015.4]
  wire [15:0] _T_21714; // @[Mux.scala 19:72:@20016.4]
  wire [7:0] _T_22292; // @[Mux.scala 19:72:@20366.4]
  wire [7:0] _T_22299; // @[Mux.scala 19:72:@20373.4]
  wire [15:0] _T_22300; // @[Mux.scala 19:72:@20374.4]
  wire [15:0] _T_22302; // @[Mux.scala 19:72:@20375.4]
  wire [7:0] _T_22309; // @[Mux.scala 19:72:@20382.4]
  wire [7:0] _T_22316; // @[Mux.scala 19:72:@20389.4]
  wire [15:0] _T_22317; // @[Mux.scala 19:72:@20390.4]
  wire [15:0] _T_22319; // @[Mux.scala 19:72:@20391.4]
  wire [7:0] _T_22326; // @[Mux.scala 19:72:@20398.4]
  wire [7:0] _T_22333; // @[Mux.scala 19:72:@20405.4]
  wire [15:0] _T_22334; // @[Mux.scala 19:72:@20406.4]
  wire [15:0] _T_22336; // @[Mux.scala 19:72:@20407.4]
  wire [7:0] _T_22343; // @[Mux.scala 19:72:@20414.4]
  wire [7:0] _T_22350; // @[Mux.scala 19:72:@20421.4]
  wire [15:0] _T_22351; // @[Mux.scala 19:72:@20422.4]
  wire [15:0] _T_22353; // @[Mux.scala 19:72:@20423.4]
  wire [7:0] _T_22360; // @[Mux.scala 19:72:@20430.4]
  wire [7:0] _T_22367; // @[Mux.scala 19:72:@20437.4]
  wire [15:0] _T_22368; // @[Mux.scala 19:72:@20438.4]
  wire [15:0] _T_22370; // @[Mux.scala 19:72:@20439.4]
  wire [7:0] _T_22377; // @[Mux.scala 19:72:@20446.4]
  wire [7:0] _T_22384; // @[Mux.scala 19:72:@20453.4]
  wire [15:0] _T_22385; // @[Mux.scala 19:72:@20454.4]
  wire [15:0] _T_22387; // @[Mux.scala 19:72:@20455.4]
  wire [7:0] _T_22394; // @[Mux.scala 19:72:@20462.4]
  wire [7:0] _T_22401; // @[Mux.scala 19:72:@20469.4]
  wire [15:0] _T_22402; // @[Mux.scala 19:72:@20470.4]
  wire [15:0] _T_22404; // @[Mux.scala 19:72:@20471.4]
  wire [7:0] _T_22411; // @[Mux.scala 19:72:@20478.4]
  wire [7:0] _T_22418; // @[Mux.scala 19:72:@20485.4]
  wire [15:0] _T_22419; // @[Mux.scala 19:72:@20486.4]
  wire [15:0] _T_22421; // @[Mux.scala 19:72:@20487.4]
  wire [15:0] _T_22436; // @[Mux.scala 19:72:@20502.4]
  wire [15:0] _T_22438; // @[Mux.scala 19:72:@20503.4]
  wire [15:0] _T_22453; // @[Mux.scala 19:72:@20518.4]
  wire [15:0] _T_22455; // @[Mux.scala 19:72:@20519.4]
  wire [15:0] _T_22470; // @[Mux.scala 19:72:@20534.4]
  wire [15:0] _T_22472; // @[Mux.scala 19:72:@20535.4]
  wire [15:0] _T_22487; // @[Mux.scala 19:72:@20550.4]
  wire [15:0] _T_22489; // @[Mux.scala 19:72:@20551.4]
  wire [15:0] _T_22504; // @[Mux.scala 19:72:@20566.4]
  wire [15:0] _T_22506; // @[Mux.scala 19:72:@20567.4]
  wire [15:0] _T_22521; // @[Mux.scala 19:72:@20582.4]
  wire [15:0] _T_22523; // @[Mux.scala 19:72:@20583.4]
  wire [15:0] _T_22538; // @[Mux.scala 19:72:@20598.4]
  wire [15:0] _T_22540; // @[Mux.scala 19:72:@20599.4]
  wire [15:0] _T_22555; // @[Mux.scala 19:72:@20614.4]
  wire [15:0] _T_22557; // @[Mux.scala 19:72:@20615.4]
  wire [15:0] _T_22558; // @[Mux.scala 19:72:@20616.4]
  wire [15:0] _T_22559; // @[Mux.scala 19:72:@20617.4]
  wire [15:0] _T_22560; // @[Mux.scala 19:72:@20618.4]
  wire [15:0] _T_22561; // @[Mux.scala 19:72:@20619.4]
  wire [15:0] _T_22562; // @[Mux.scala 19:72:@20620.4]
  wire [15:0] _T_22563; // @[Mux.scala 19:72:@20621.4]
  wire [15:0] _T_22564; // @[Mux.scala 19:72:@20622.4]
  wire [15:0] _T_22565; // @[Mux.scala 19:72:@20623.4]
  wire [15:0] _T_22566; // @[Mux.scala 19:72:@20624.4]
  wire [15:0] _T_22567; // @[Mux.scala 19:72:@20625.4]
  wire [15:0] _T_22568; // @[Mux.scala 19:72:@20626.4]
  wire [15:0] _T_22569; // @[Mux.scala 19:72:@20627.4]
  wire [15:0] _T_22570; // @[Mux.scala 19:72:@20628.4]
  wire [15:0] _T_22571; // @[Mux.scala 19:72:@20629.4]
  wire [15:0] _T_22572; // @[Mux.scala 19:72:@20630.4]
  wire [7:0] _T_23150; // @[Mux.scala 19:72:@20980.4]
  wire [7:0] _T_23157; // @[Mux.scala 19:72:@20987.4]
  wire [15:0] _T_23158; // @[Mux.scala 19:72:@20988.4]
  wire [15:0] _T_23160; // @[Mux.scala 19:72:@20989.4]
  wire [7:0] _T_23167; // @[Mux.scala 19:72:@20996.4]
  wire [7:0] _T_23174; // @[Mux.scala 19:72:@21003.4]
  wire [15:0] _T_23175; // @[Mux.scala 19:72:@21004.4]
  wire [15:0] _T_23177; // @[Mux.scala 19:72:@21005.4]
  wire [7:0] _T_23184; // @[Mux.scala 19:72:@21012.4]
  wire [7:0] _T_23191; // @[Mux.scala 19:72:@21019.4]
  wire [15:0] _T_23192; // @[Mux.scala 19:72:@21020.4]
  wire [15:0] _T_23194; // @[Mux.scala 19:72:@21021.4]
  wire [7:0] _T_23201; // @[Mux.scala 19:72:@21028.4]
  wire [7:0] _T_23208; // @[Mux.scala 19:72:@21035.4]
  wire [15:0] _T_23209; // @[Mux.scala 19:72:@21036.4]
  wire [15:0] _T_23211; // @[Mux.scala 19:72:@21037.4]
  wire [7:0] _T_23218; // @[Mux.scala 19:72:@21044.4]
  wire [7:0] _T_23225; // @[Mux.scala 19:72:@21051.4]
  wire [15:0] _T_23226; // @[Mux.scala 19:72:@21052.4]
  wire [15:0] _T_23228; // @[Mux.scala 19:72:@21053.4]
  wire [7:0] _T_23235; // @[Mux.scala 19:72:@21060.4]
  wire [7:0] _T_23242; // @[Mux.scala 19:72:@21067.4]
  wire [15:0] _T_23243; // @[Mux.scala 19:72:@21068.4]
  wire [15:0] _T_23245; // @[Mux.scala 19:72:@21069.4]
  wire [7:0] _T_23252; // @[Mux.scala 19:72:@21076.4]
  wire [7:0] _T_23259; // @[Mux.scala 19:72:@21083.4]
  wire [15:0] _T_23260; // @[Mux.scala 19:72:@21084.4]
  wire [15:0] _T_23262; // @[Mux.scala 19:72:@21085.4]
  wire [7:0] _T_23269; // @[Mux.scala 19:72:@21092.4]
  wire [7:0] _T_23276; // @[Mux.scala 19:72:@21099.4]
  wire [15:0] _T_23277; // @[Mux.scala 19:72:@21100.4]
  wire [15:0] _T_23279; // @[Mux.scala 19:72:@21101.4]
  wire [15:0] _T_23294; // @[Mux.scala 19:72:@21116.4]
  wire [15:0] _T_23296; // @[Mux.scala 19:72:@21117.4]
  wire [15:0] _T_23311; // @[Mux.scala 19:72:@21132.4]
  wire [15:0] _T_23313; // @[Mux.scala 19:72:@21133.4]
  wire [15:0] _T_23328; // @[Mux.scala 19:72:@21148.4]
  wire [15:0] _T_23330; // @[Mux.scala 19:72:@21149.4]
  wire [15:0] _T_23345; // @[Mux.scala 19:72:@21164.4]
  wire [15:0] _T_23347; // @[Mux.scala 19:72:@21165.4]
  wire [15:0] _T_23362; // @[Mux.scala 19:72:@21180.4]
  wire [15:0] _T_23364; // @[Mux.scala 19:72:@21181.4]
  wire [15:0] _T_23379; // @[Mux.scala 19:72:@21196.4]
  wire [15:0] _T_23381; // @[Mux.scala 19:72:@21197.4]
  wire [15:0] _T_23396; // @[Mux.scala 19:72:@21212.4]
  wire [15:0] _T_23398; // @[Mux.scala 19:72:@21213.4]
  wire [15:0] _T_23413; // @[Mux.scala 19:72:@21228.4]
  wire [15:0] _T_23415; // @[Mux.scala 19:72:@21229.4]
  wire [15:0] _T_23416; // @[Mux.scala 19:72:@21230.4]
  wire [15:0] _T_23417; // @[Mux.scala 19:72:@21231.4]
  wire [15:0] _T_23418; // @[Mux.scala 19:72:@21232.4]
  wire [15:0] _T_23419; // @[Mux.scala 19:72:@21233.4]
  wire [15:0] _T_23420; // @[Mux.scala 19:72:@21234.4]
  wire [15:0] _T_23421; // @[Mux.scala 19:72:@21235.4]
  wire [15:0] _T_23422; // @[Mux.scala 19:72:@21236.4]
  wire [15:0] _T_23423; // @[Mux.scala 19:72:@21237.4]
  wire [15:0] _T_23424; // @[Mux.scala 19:72:@21238.4]
  wire [15:0] _T_23425; // @[Mux.scala 19:72:@21239.4]
  wire [15:0] _T_23426; // @[Mux.scala 19:72:@21240.4]
  wire [15:0] _T_23427; // @[Mux.scala 19:72:@21241.4]
  wire [15:0] _T_23428; // @[Mux.scala 19:72:@21242.4]
  wire [15:0] _T_23429; // @[Mux.scala 19:72:@21243.4]
  wire [15:0] _T_23430; // @[Mux.scala 19:72:@21244.4]
  wire [7:0] _T_24008; // @[Mux.scala 19:72:@21594.4]
  wire [7:0] _T_24015; // @[Mux.scala 19:72:@21601.4]
  wire [15:0] _T_24016; // @[Mux.scala 19:72:@21602.4]
  wire [15:0] _T_24018; // @[Mux.scala 19:72:@21603.4]
  wire [7:0] _T_24025; // @[Mux.scala 19:72:@21610.4]
  wire [7:0] _T_24032; // @[Mux.scala 19:72:@21617.4]
  wire [15:0] _T_24033; // @[Mux.scala 19:72:@21618.4]
  wire [15:0] _T_24035; // @[Mux.scala 19:72:@21619.4]
  wire [7:0] _T_24042; // @[Mux.scala 19:72:@21626.4]
  wire [7:0] _T_24049; // @[Mux.scala 19:72:@21633.4]
  wire [15:0] _T_24050; // @[Mux.scala 19:72:@21634.4]
  wire [15:0] _T_24052; // @[Mux.scala 19:72:@21635.4]
  wire [7:0] _T_24059; // @[Mux.scala 19:72:@21642.4]
  wire [7:0] _T_24066; // @[Mux.scala 19:72:@21649.4]
  wire [15:0] _T_24067; // @[Mux.scala 19:72:@21650.4]
  wire [15:0] _T_24069; // @[Mux.scala 19:72:@21651.4]
  wire [7:0] _T_24076; // @[Mux.scala 19:72:@21658.4]
  wire [7:0] _T_24083; // @[Mux.scala 19:72:@21665.4]
  wire [15:0] _T_24084; // @[Mux.scala 19:72:@21666.4]
  wire [15:0] _T_24086; // @[Mux.scala 19:72:@21667.4]
  wire [7:0] _T_24093; // @[Mux.scala 19:72:@21674.4]
  wire [7:0] _T_24100; // @[Mux.scala 19:72:@21681.4]
  wire [15:0] _T_24101; // @[Mux.scala 19:72:@21682.4]
  wire [15:0] _T_24103; // @[Mux.scala 19:72:@21683.4]
  wire [7:0] _T_24110; // @[Mux.scala 19:72:@21690.4]
  wire [7:0] _T_24117; // @[Mux.scala 19:72:@21697.4]
  wire [15:0] _T_24118; // @[Mux.scala 19:72:@21698.4]
  wire [15:0] _T_24120; // @[Mux.scala 19:72:@21699.4]
  wire [7:0] _T_24127; // @[Mux.scala 19:72:@21706.4]
  wire [7:0] _T_24134; // @[Mux.scala 19:72:@21713.4]
  wire [15:0] _T_24135; // @[Mux.scala 19:72:@21714.4]
  wire [15:0] _T_24137; // @[Mux.scala 19:72:@21715.4]
  wire [15:0] _T_24152; // @[Mux.scala 19:72:@21730.4]
  wire [15:0] _T_24154; // @[Mux.scala 19:72:@21731.4]
  wire [15:0] _T_24169; // @[Mux.scala 19:72:@21746.4]
  wire [15:0] _T_24171; // @[Mux.scala 19:72:@21747.4]
  wire [15:0] _T_24186; // @[Mux.scala 19:72:@21762.4]
  wire [15:0] _T_24188; // @[Mux.scala 19:72:@21763.4]
  wire [15:0] _T_24203; // @[Mux.scala 19:72:@21778.4]
  wire [15:0] _T_24205; // @[Mux.scala 19:72:@21779.4]
  wire [15:0] _T_24220; // @[Mux.scala 19:72:@21794.4]
  wire [15:0] _T_24222; // @[Mux.scala 19:72:@21795.4]
  wire [15:0] _T_24237; // @[Mux.scala 19:72:@21810.4]
  wire [15:0] _T_24239; // @[Mux.scala 19:72:@21811.4]
  wire [15:0] _T_24254; // @[Mux.scala 19:72:@21826.4]
  wire [15:0] _T_24256; // @[Mux.scala 19:72:@21827.4]
  wire [15:0] _T_24271; // @[Mux.scala 19:72:@21842.4]
  wire [15:0] _T_24273; // @[Mux.scala 19:72:@21843.4]
  wire [15:0] _T_24274; // @[Mux.scala 19:72:@21844.4]
  wire [15:0] _T_24275; // @[Mux.scala 19:72:@21845.4]
  wire [15:0] _T_24276; // @[Mux.scala 19:72:@21846.4]
  wire [15:0] _T_24277; // @[Mux.scala 19:72:@21847.4]
  wire [15:0] _T_24278; // @[Mux.scala 19:72:@21848.4]
  wire [15:0] _T_24279; // @[Mux.scala 19:72:@21849.4]
  wire [15:0] _T_24280; // @[Mux.scala 19:72:@21850.4]
  wire [15:0] _T_24281; // @[Mux.scala 19:72:@21851.4]
  wire [15:0] _T_24282; // @[Mux.scala 19:72:@21852.4]
  wire [15:0] _T_24283; // @[Mux.scala 19:72:@21853.4]
  wire [15:0] _T_24284; // @[Mux.scala 19:72:@21854.4]
  wire [15:0] _T_24285; // @[Mux.scala 19:72:@21855.4]
  wire [15:0] _T_24286; // @[Mux.scala 19:72:@21856.4]
  wire [15:0] _T_24287; // @[Mux.scala 19:72:@21857.4]
  wire [15:0] _T_24288; // @[Mux.scala 19:72:@21858.4]
  wire [7:0] _T_24866; // @[Mux.scala 19:72:@22208.4]
  wire [7:0] _T_24873; // @[Mux.scala 19:72:@22215.4]
  wire [15:0] _T_24874; // @[Mux.scala 19:72:@22216.4]
  wire [15:0] _T_24876; // @[Mux.scala 19:72:@22217.4]
  wire [7:0] _T_24883; // @[Mux.scala 19:72:@22224.4]
  wire [7:0] _T_24890; // @[Mux.scala 19:72:@22231.4]
  wire [15:0] _T_24891; // @[Mux.scala 19:72:@22232.4]
  wire [15:0] _T_24893; // @[Mux.scala 19:72:@22233.4]
  wire [7:0] _T_24900; // @[Mux.scala 19:72:@22240.4]
  wire [7:0] _T_24907; // @[Mux.scala 19:72:@22247.4]
  wire [15:0] _T_24908; // @[Mux.scala 19:72:@22248.4]
  wire [15:0] _T_24910; // @[Mux.scala 19:72:@22249.4]
  wire [7:0] _T_24917; // @[Mux.scala 19:72:@22256.4]
  wire [7:0] _T_24924; // @[Mux.scala 19:72:@22263.4]
  wire [15:0] _T_24925; // @[Mux.scala 19:72:@22264.4]
  wire [15:0] _T_24927; // @[Mux.scala 19:72:@22265.4]
  wire [7:0] _T_24934; // @[Mux.scala 19:72:@22272.4]
  wire [7:0] _T_24941; // @[Mux.scala 19:72:@22279.4]
  wire [15:0] _T_24942; // @[Mux.scala 19:72:@22280.4]
  wire [15:0] _T_24944; // @[Mux.scala 19:72:@22281.4]
  wire [7:0] _T_24951; // @[Mux.scala 19:72:@22288.4]
  wire [7:0] _T_24958; // @[Mux.scala 19:72:@22295.4]
  wire [15:0] _T_24959; // @[Mux.scala 19:72:@22296.4]
  wire [15:0] _T_24961; // @[Mux.scala 19:72:@22297.4]
  wire [7:0] _T_24968; // @[Mux.scala 19:72:@22304.4]
  wire [7:0] _T_24975; // @[Mux.scala 19:72:@22311.4]
  wire [15:0] _T_24976; // @[Mux.scala 19:72:@22312.4]
  wire [15:0] _T_24978; // @[Mux.scala 19:72:@22313.4]
  wire [7:0] _T_24985; // @[Mux.scala 19:72:@22320.4]
  wire [7:0] _T_24992; // @[Mux.scala 19:72:@22327.4]
  wire [15:0] _T_24993; // @[Mux.scala 19:72:@22328.4]
  wire [15:0] _T_24995; // @[Mux.scala 19:72:@22329.4]
  wire [15:0] _T_25010; // @[Mux.scala 19:72:@22344.4]
  wire [15:0] _T_25012; // @[Mux.scala 19:72:@22345.4]
  wire [15:0] _T_25027; // @[Mux.scala 19:72:@22360.4]
  wire [15:0] _T_25029; // @[Mux.scala 19:72:@22361.4]
  wire [15:0] _T_25044; // @[Mux.scala 19:72:@22376.4]
  wire [15:0] _T_25046; // @[Mux.scala 19:72:@22377.4]
  wire [15:0] _T_25061; // @[Mux.scala 19:72:@22392.4]
  wire [15:0] _T_25063; // @[Mux.scala 19:72:@22393.4]
  wire [15:0] _T_25078; // @[Mux.scala 19:72:@22408.4]
  wire [15:0] _T_25080; // @[Mux.scala 19:72:@22409.4]
  wire [15:0] _T_25095; // @[Mux.scala 19:72:@22424.4]
  wire [15:0] _T_25097; // @[Mux.scala 19:72:@22425.4]
  wire [15:0] _T_25112; // @[Mux.scala 19:72:@22440.4]
  wire [15:0] _T_25114; // @[Mux.scala 19:72:@22441.4]
  wire [15:0] _T_25129; // @[Mux.scala 19:72:@22456.4]
  wire [15:0] _T_25131; // @[Mux.scala 19:72:@22457.4]
  wire [15:0] _T_25132; // @[Mux.scala 19:72:@22458.4]
  wire [15:0] _T_25133; // @[Mux.scala 19:72:@22459.4]
  wire [15:0] _T_25134; // @[Mux.scala 19:72:@22460.4]
  wire [15:0] _T_25135; // @[Mux.scala 19:72:@22461.4]
  wire [15:0] _T_25136; // @[Mux.scala 19:72:@22462.4]
  wire [15:0] _T_25137; // @[Mux.scala 19:72:@22463.4]
  wire [15:0] _T_25138; // @[Mux.scala 19:72:@22464.4]
  wire [15:0] _T_25139; // @[Mux.scala 19:72:@22465.4]
  wire [15:0] _T_25140; // @[Mux.scala 19:72:@22466.4]
  wire [15:0] _T_25141; // @[Mux.scala 19:72:@22467.4]
  wire [15:0] _T_25142; // @[Mux.scala 19:72:@22468.4]
  wire [15:0] _T_25143; // @[Mux.scala 19:72:@22469.4]
  wire [15:0] _T_25144; // @[Mux.scala 19:72:@22470.4]
  wire [15:0] _T_25145; // @[Mux.scala 19:72:@22471.4]
  wire [15:0] _T_25146; // @[Mux.scala 19:72:@22472.4]
  wire [7:0] _T_25724; // @[Mux.scala 19:72:@22822.4]
  wire [7:0] _T_25731; // @[Mux.scala 19:72:@22829.4]
  wire [15:0] _T_25732; // @[Mux.scala 19:72:@22830.4]
  wire [15:0] _T_25734; // @[Mux.scala 19:72:@22831.4]
  wire [7:0] _T_25741; // @[Mux.scala 19:72:@22838.4]
  wire [7:0] _T_25748; // @[Mux.scala 19:72:@22845.4]
  wire [15:0] _T_25749; // @[Mux.scala 19:72:@22846.4]
  wire [15:0] _T_25751; // @[Mux.scala 19:72:@22847.4]
  wire [7:0] _T_25758; // @[Mux.scala 19:72:@22854.4]
  wire [7:0] _T_25765; // @[Mux.scala 19:72:@22861.4]
  wire [15:0] _T_25766; // @[Mux.scala 19:72:@22862.4]
  wire [15:0] _T_25768; // @[Mux.scala 19:72:@22863.4]
  wire [7:0] _T_25775; // @[Mux.scala 19:72:@22870.4]
  wire [7:0] _T_25782; // @[Mux.scala 19:72:@22877.4]
  wire [15:0] _T_25783; // @[Mux.scala 19:72:@22878.4]
  wire [15:0] _T_25785; // @[Mux.scala 19:72:@22879.4]
  wire [7:0] _T_25792; // @[Mux.scala 19:72:@22886.4]
  wire [7:0] _T_25799; // @[Mux.scala 19:72:@22893.4]
  wire [15:0] _T_25800; // @[Mux.scala 19:72:@22894.4]
  wire [15:0] _T_25802; // @[Mux.scala 19:72:@22895.4]
  wire [7:0] _T_25809; // @[Mux.scala 19:72:@22902.4]
  wire [7:0] _T_25816; // @[Mux.scala 19:72:@22909.4]
  wire [15:0] _T_25817; // @[Mux.scala 19:72:@22910.4]
  wire [15:0] _T_25819; // @[Mux.scala 19:72:@22911.4]
  wire [7:0] _T_25826; // @[Mux.scala 19:72:@22918.4]
  wire [7:0] _T_25833; // @[Mux.scala 19:72:@22925.4]
  wire [15:0] _T_25834; // @[Mux.scala 19:72:@22926.4]
  wire [15:0] _T_25836; // @[Mux.scala 19:72:@22927.4]
  wire [7:0] _T_25843; // @[Mux.scala 19:72:@22934.4]
  wire [7:0] _T_25850; // @[Mux.scala 19:72:@22941.4]
  wire [15:0] _T_25851; // @[Mux.scala 19:72:@22942.4]
  wire [15:0] _T_25853; // @[Mux.scala 19:72:@22943.4]
  wire [15:0] _T_25868; // @[Mux.scala 19:72:@22958.4]
  wire [15:0] _T_25870; // @[Mux.scala 19:72:@22959.4]
  wire [15:0] _T_25885; // @[Mux.scala 19:72:@22974.4]
  wire [15:0] _T_25887; // @[Mux.scala 19:72:@22975.4]
  wire [15:0] _T_25902; // @[Mux.scala 19:72:@22990.4]
  wire [15:0] _T_25904; // @[Mux.scala 19:72:@22991.4]
  wire [15:0] _T_25919; // @[Mux.scala 19:72:@23006.4]
  wire [15:0] _T_25921; // @[Mux.scala 19:72:@23007.4]
  wire [15:0] _T_25936; // @[Mux.scala 19:72:@23022.4]
  wire [15:0] _T_25938; // @[Mux.scala 19:72:@23023.4]
  wire [15:0] _T_25953; // @[Mux.scala 19:72:@23038.4]
  wire [15:0] _T_25955; // @[Mux.scala 19:72:@23039.4]
  wire [15:0] _T_25970; // @[Mux.scala 19:72:@23054.4]
  wire [15:0] _T_25972; // @[Mux.scala 19:72:@23055.4]
  wire [15:0] _T_25987; // @[Mux.scala 19:72:@23070.4]
  wire [15:0] _T_25989; // @[Mux.scala 19:72:@23071.4]
  wire [15:0] _T_25990; // @[Mux.scala 19:72:@23072.4]
  wire [15:0] _T_25991; // @[Mux.scala 19:72:@23073.4]
  wire [15:0] _T_25992; // @[Mux.scala 19:72:@23074.4]
  wire [15:0] _T_25993; // @[Mux.scala 19:72:@23075.4]
  wire [15:0] _T_25994; // @[Mux.scala 19:72:@23076.4]
  wire [15:0] _T_25995; // @[Mux.scala 19:72:@23077.4]
  wire [15:0] _T_25996; // @[Mux.scala 19:72:@23078.4]
  wire [15:0] _T_25997; // @[Mux.scala 19:72:@23079.4]
  wire [15:0] _T_25998; // @[Mux.scala 19:72:@23080.4]
  wire [15:0] _T_25999; // @[Mux.scala 19:72:@23081.4]
  wire [15:0] _T_26000; // @[Mux.scala 19:72:@23082.4]
  wire [15:0] _T_26001; // @[Mux.scala 19:72:@23083.4]
  wire [15:0] _T_26002; // @[Mux.scala 19:72:@23084.4]
  wire [15:0] _T_26003; // @[Mux.scala 19:72:@23085.4]
  wire [15:0] _T_26004; // @[Mux.scala 19:72:@23086.4]
  wire [7:0] _T_26582; // @[Mux.scala 19:72:@23436.4]
  wire [7:0] _T_26589; // @[Mux.scala 19:72:@23443.4]
  wire [15:0] _T_26590; // @[Mux.scala 19:72:@23444.4]
  wire [15:0] _T_26592; // @[Mux.scala 19:72:@23445.4]
  wire [7:0] _T_26599; // @[Mux.scala 19:72:@23452.4]
  wire [7:0] _T_26606; // @[Mux.scala 19:72:@23459.4]
  wire [15:0] _T_26607; // @[Mux.scala 19:72:@23460.4]
  wire [15:0] _T_26609; // @[Mux.scala 19:72:@23461.4]
  wire [7:0] _T_26616; // @[Mux.scala 19:72:@23468.4]
  wire [7:0] _T_26623; // @[Mux.scala 19:72:@23475.4]
  wire [15:0] _T_26624; // @[Mux.scala 19:72:@23476.4]
  wire [15:0] _T_26626; // @[Mux.scala 19:72:@23477.4]
  wire [7:0] _T_26633; // @[Mux.scala 19:72:@23484.4]
  wire [7:0] _T_26640; // @[Mux.scala 19:72:@23491.4]
  wire [15:0] _T_26641; // @[Mux.scala 19:72:@23492.4]
  wire [15:0] _T_26643; // @[Mux.scala 19:72:@23493.4]
  wire [7:0] _T_26650; // @[Mux.scala 19:72:@23500.4]
  wire [7:0] _T_26657; // @[Mux.scala 19:72:@23507.4]
  wire [15:0] _T_26658; // @[Mux.scala 19:72:@23508.4]
  wire [15:0] _T_26660; // @[Mux.scala 19:72:@23509.4]
  wire [7:0] _T_26667; // @[Mux.scala 19:72:@23516.4]
  wire [7:0] _T_26674; // @[Mux.scala 19:72:@23523.4]
  wire [15:0] _T_26675; // @[Mux.scala 19:72:@23524.4]
  wire [15:0] _T_26677; // @[Mux.scala 19:72:@23525.4]
  wire [7:0] _T_26684; // @[Mux.scala 19:72:@23532.4]
  wire [7:0] _T_26691; // @[Mux.scala 19:72:@23539.4]
  wire [15:0] _T_26692; // @[Mux.scala 19:72:@23540.4]
  wire [15:0] _T_26694; // @[Mux.scala 19:72:@23541.4]
  wire [7:0] _T_26701; // @[Mux.scala 19:72:@23548.4]
  wire [7:0] _T_26708; // @[Mux.scala 19:72:@23555.4]
  wire [15:0] _T_26709; // @[Mux.scala 19:72:@23556.4]
  wire [15:0] _T_26711; // @[Mux.scala 19:72:@23557.4]
  wire [15:0] _T_26726; // @[Mux.scala 19:72:@23572.4]
  wire [15:0] _T_26728; // @[Mux.scala 19:72:@23573.4]
  wire [15:0] _T_26743; // @[Mux.scala 19:72:@23588.4]
  wire [15:0] _T_26745; // @[Mux.scala 19:72:@23589.4]
  wire [15:0] _T_26760; // @[Mux.scala 19:72:@23604.4]
  wire [15:0] _T_26762; // @[Mux.scala 19:72:@23605.4]
  wire [15:0] _T_26777; // @[Mux.scala 19:72:@23620.4]
  wire [15:0] _T_26779; // @[Mux.scala 19:72:@23621.4]
  wire [15:0] _T_26794; // @[Mux.scala 19:72:@23636.4]
  wire [15:0] _T_26796; // @[Mux.scala 19:72:@23637.4]
  wire [15:0] _T_26811; // @[Mux.scala 19:72:@23652.4]
  wire [15:0] _T_26813; // @[Mux.scala 19:72:@23653.4]
  wire [15:0] _T_26828; // @[Mux.scala 19:72:@23668.4]
  wire [15:0] _T_26830; // @[Mux.scala 19:72:@23669.4]
  wire [15:0] _T_26845; // @[Mux.scala 19:72:@23684.4]
  wire [15:0] _T_26847; // @[Mux.scala 19:72:@23685.4]
  wire [15:0] _T_26848; // @[Mux.scala 19:72:@23686.4]
  wire [15:0] _T_26849; // @[Mux.scala 19:72:@23687.4]
  wire [15:0] _T_26850; // @[Mux.scala 19:72:@23688.4]
  wire [15:0] _T_26851; // @[Mux.scala 19:72:@23689.4]
  wire [15:0] _T_26852; // @[Mux.scala 19:72:@23690.4]
  wire [15:0] _T_26853; // @[Mux.scala 19:72:@23691.4]
  wire [15:0] _T_26854; // @[Mux.scala 19:72:@23692.4]
  wire [15:0] _T_26855; // @[Mux.scala 19:72:@23693.4]
  wire [15:0] _T_26856; // @[Mux.scala 19:72:@23694.4]
  wire [15:0] _T_26857; // @[Mux.scala 19:72:@23695.4]
  wire [15:0] _T_26858; // @[Mux.scala 19:72:@23696.4]
  wire [15:0] _T_26859; // @[Mux.scala 19:72:@23697.4]
  wire [15:0] _T_26860; // @[Mux.scala 19:72:@23698.4]
  wire [15:0] _T_26861; // @[Mux.scala 19:72:@23699.4]
  wire [15:0] _T_26862; // @[Mux.scala 19:72:@23700.4]
  wire [7:0] _T_27440; // @[Mux.scala 19:72:@24050.4]
  wire [7:0] _T_27447; // @[Mux.scala 19:72:@24057.4]
  wire [15:0] _T_27448; // @[Mux.scala 19:72:@24058.4]
  wire [15:0] _T_27450; // @[Mux.scala 19:72:@24059.4]
  wire [7:0] _T_27457; // @[Mux.scala 19:72:@24066.4]
  wire [7:0] _T_27464; // @[Mux.scala 19:72:@24073.4]
  wire [15:0] _T_27465; // @[Mux.scala 19:72:@24074.4]
  wire [15:0] _T_27467; // @[Mux.scala 19:72:@24075.4]
  wire [7:0] _T_27474; // @[Mux.scala 19:72:@24082.4]
  wire [7:0] _T_27481; // @[Mux.scala 19:72:@24089.4]
  wire [15:0] _T_27482; // @[Mux.scala 19:72:@24090.4]
  wire [15:0] _T_27484; // @[Mux.scala 19:72:@24091.4]
  wire [7:0] _T_27491; // @[Mux.scala 19:72:@24098.4]
  wire [7:0] _T_27498; // @[Mux.scala 19:72:@24105.4]
  wire [15:0] _T_27499; // @[Mux.scala 19:72:@24106.4]
  wire [15:0] _T_27501; // @[Mux.scala 19:72:@24107.4]
  wire [7:0] _T_27508; // @[Mux.scala 19:72:@24114.4]
  wire [7:0] _T_27515; // @[Mux.scala 19:72:@24121.4]
  wire [15:0] _T_27516; // @[Mux.scala 19:72:@24122.4]
  wire [15:0] _T_27518; // @[Mux.scala 19:72:@24123.4]
  wire [7:0] _T_27525; // @[Mux.scala 19:72:@24130.4]
  wire [7:0] _T_27532; // @[Mux.scala 19:72:@24137.4]
  wire [15:0] _T_27533; // @[Mux.scala 19:72:@24138.4]
  wire [15:0] _T_27535; // @[Mux.scala 19:72:@24139.4]
  wire [7:0] _T_27542; // @[Mux.scala 19:72:@24146.4]
  wire [7:0] _T_27549; // @[Mux.scala 19:72:@24153.4]
  wire [15:0] _T_27550; // @[Mux.scala 19:72:@24154.4]
  wire [15:0] _T_27552; // @[Mux.scala 19:72:@24155.4]
  wire [7:0] _T_27559; // @[Mux.scala 19:72:@24162.4]
  wire [7:0] _T_27566; // @[Mux.scala 19:72:@24169.4]
  wire [15:0] _T_27567; // @[Mux.scala 19:72:@24170.4]
  wire [15:0] _T_27569; // @[Mux.scala 19:72:@24171.4]
  wire [15:0] _T_27584; // @[Mux.scala 19:72:@24186.4]
  wire [15:0] _T_27586; // @[Mux.scala 19:72:@24187.4]
  wire [15:0] _T_27601; // @[Mux.scala 19:72:@24202.4]
  wire [15:0] _T_27603; // @[Mux.scala 19:72:@24203.4]
  wire [15:0] _T_27618; // @[Mux.scala 19:72:@24218.4]
  wire [15:0] _T_27620; // @[Mux.scala 19:72:@24219.4]
  wire [15:0] _T_27635; // @[Mux.scala 19:72:@24234.4]
  wire [15:0] _T_27637; // @[Mux.scala 19:72:@24235.4]
  wire [15:0] _T_27652; // @[Mux.scala 19:72:@24250.4]
  wire [15:0] _T_27654; // @[Mux.scala 19:72:@24251.4]
  wire [15:0] _T_27669; // @[Mux.scala 19:72:@24266.4]
  wire [15:0] _T_27671; // @[Mux.scala 19:72:@24267.4]
  wire [15:0] _T_27686; // @[Mux.scala 19:72:@24282.4]
  wire [15:0] _T_27688; // @[Mux.scala 19:72:@24283.4]
  wire [15:0] _T_27703; // @[Mux.scala 19:72:@24298.4]
  wire [15:0] _T_27705; // @[Mux.scala 19:72:@24299.4]
  wire [15:0] _T_27706; // @[Mux.scala 19:72:@24300.4]
  wire [15:0] _T_27707; // @[Mux.scala 19:72:@24301.4]
  wire [15:0] _T_27708; // @[Mux.scala 19:72:@24302.4]
  wire [15:0] _T_27709; // @[Mux.scala 19:72:@24303.4]
  wire [15:0] _T_27710; // @[Mux.scala 19:72:@24304.4]
  wire [15:0] _T_27711; // @[Mux.scala 19:72:@24305.4]
  wire [15:0] _T_27712; // @[Mux.scala 19:72:@24306.4]
  wire [15:0] _T_27713; // @[Mux.scala 19:72:@24307.4]
  wire [15:0] _T_27714; // @[Mux.scala 19:72:@24308.4]
  wire [15:0] _T_27715; // @[Mux.scala 19:72:@24309.4]
  wire [15:0] _T_27716; // @[Mux.scala 19:72:@24310.4]
  wire [15:0] _T_27717; // @[Mux.scala 19:72:@24311.4]
  wire [15:0] _T_27718; // @[Mux.scala 19:72:@24312.4]
  wire [15:0] _T_27719; // @[Mux.scala 19:72:@24313.4]
  wire [15:0] _T_27720; // @[Mux.scala 19:72:@24314.4]
  wire [7:0] _T_28298; // @[Mux.scala 19:72:@24664.4]
  wire [7:0] _T_28305; // @[Mux.scala 19:72:@24671.4]
  wire [15:0] _T_28306; // @[Mux.scala 19:72:@24672.4]
  wire [15:0] _T_28308; // @[Mux.scala 19:72:@24673.4]
  wire [7:0] _T_28315; // @[Mux.scala 19:72:@24680.4]
  wire [7:0] _T_28322; // @[Mux.scala 19:72:@24687.4]
  wire [15:0] _T_28323; // @[Mux.scala 19:72:@24688.4]
  wire [15:0] _T_28325; // @[Mux.scala 19:72:@24689.4]
  wire [7:0] _T_28332; // @[Mux.scala 19:72:@24696.4]
  wire [7:0] _T_28339; // @[Mux.scala 19:72:@24703.4]
  wire [15:0] _T_28340; // @[Mux.scala 19:72:@24704.4]
  wire [15:0] _T_28342; // @[Mux.scala 19:72:@24705.4]
  wire [7:0] _T_28349; // @[Mux.scala 19:72:@24712.4]
  wire [7:0] _T_28356; // @[Mux.scala 19:72:@24719.4]
  wire [15:0] _T_28357; // @[Mux.scala 19:72:@24720.4]
  wire [15:0] _T_28359; // @[Mux.scala 19:72:@24721.4]
  wire [7:0] _T_28366; // @[Mux.scala 19:72:@24728.4]
  wire [7:0] _T_28373; // @[Mux.scala 19:72:@24735.4]
  wire [15:0] _T_28374; // @[Mux.scala 19:72:@24736.4]
  wire [15:0] _T_28376; // @[Mux.scala 19:72:@24737.4]
  wire [7:0] _T_28383; // @[Mux.scala 19:72:@24744.4]
  wire [7:0] _T_28390; // @[Mux.scala 19:72:@24751.4]
  wire [15:0] _T_28391; // @[Mux.scala 19:72:@24752.4]
  wire [15:0] _T_28393; // @[Mux.scala 19:72:@24753.4]
  wire [7:0] _T_28400; // @[Mux.scala 19:72:@24760.4]
  wire [7:0] _T_28407; // @[Mux.scala 19:72:@24767.4]
  wire [15:0] _T_28408; // @[Mux.scala 19:72:@24768.4]
  wire [15:0] _T_28410; // @[Mux.scala 19:72:@24769.4]
  wire [7:0] _T_28417; // @[Mux.scala 19:72:@24776.4]
  wire [7:0] _T_28424; // @[Mux.scala 19:72:@24783.4]
  wire [15:0] _T_28425; // @[Mux.scala 19:72:@24784.4]
  wire [15:0] _T_28427; // @[Mux.scala 19:72:@24785.4]
  wire [15:0] _T_28442; // @[Mux.scala 19:72:@24800.4]
  wire [15:0] _T_28444; // @[Mux.scala 19:72:@24801.4]
  wire [15:0] _T_28459; // @[Mux.scala 19:72:@24816.4]
  wire [15:0] _T_28461; // @[Mux.scala 19:72:@24817.4]
  wire [15:0] _T_28476; // @[Mux.scala 19:72:@24832.4]
  wire [15:0] _T_28478; // @[Mux.scala 19:72:@24833.4]
  wire [15:0] _T_28493; // @[Mux.scala 19:72:@24848.4]
  wire [15:0] _T_28495; // @[Mux.scala 19:72:@24849.4]
  wire [15:0] _T_28510; // @[Mux.scala 19:72:@24864.4]
  wire [15:0] _T_28512; // @[Mux.scala 19:72:@24865.4]
  wire [15:0] _T_28527; // @[Mux.scala 19:72:@24880.4]
  wire [15:0] _T_28529; // @[Mux.scala 19:72:@24881.4]
  wire [15:0] _T_28544; // @[Mux.scala 19:72:@24896.4]
  wire [15:0] _T_28546; // @[Mux.scala 19:72:@24897.4]
  wire [15:0] _T_28561; // @[Mux.scala 19:72:@24912.4]
  wire [15:0] _T_28563; // @[Mux.scala 19:72:@24913.4]
  wire [15:0] _T_28564; // @[Mux.scala 19:72:@24914.4]
  wire [15:0] _T_28565; // @[Mux.scala 19:72:@24915.4]
  wire [15:0] _T_28566; // @[Mux.scala 19:72:@24916.4]
  wire [15:0] _T_28567; // @[Mux.scala 19:72:@24917.4]
  wire [15:0] _T_28568; // @[Mux.scala 19:72:@24918.4]
  wire [15:0] _T_28569; // @[Mux.scala 19:72:@24919.4]
  wire [15:0] _T_28570; // @[Mux.scala 19:72:@24920.4]
  wire [15:0] _T_28571; // @[Mux.scala 19:72:@24921.4]
  wire [15:0] _T_28572; // @[Mux.scala 19:72:@24922.4]
  wire [15:0] _T_28573; // @[Mux.scala 19:72:@24923.4]
  wire [15:0] _T_28574; // @[Mux.scala 19:72:@24924.4]
  wire [15:0] _T_28575; // @[Mux.scala 19:72:@24925.4]
  wire [15:0] _T_28576; // @[Mux.scala 19:72:@24926.4]
  wire [15:0] _T_28577; // @[Mux.scala 19:72:@24927.4]
  wire [15:0] _T_28578; // @[Mux.scala 19:72:@24928.4]
  wire [7:0] _T_29156; // @[Mux.scala 19:72:@25278.4]
  wire [7:0] _T_29163; // @[Mux.scala 19:72:@25285.4]
  wire [15:0] _T_29164; // @[Mux.scala 19:72:@25286.4]
  wire [15:0] _T_29166; // @[Mux.scala 19:72:@25287.4]
  wire [7:0] _T_29173; // @[Mux.scala 19:72:@25294.4]
  wire [7:0] _T_29180; // @[Mux.scala 19:72:@25301.4]
  wire [15:0] _T_29181; // @[Mux.scala 19:72:@25302.4]
  wire [15:0] _T_29183; // @[Mux.scala 19:72:@25303.4]
  wire [7:0] _T_29190; // @[Mux.scala 19:72:@25310.4]
  wire [7:0] _T_29197; // @[Mux.scala 19:72:@25317.4]
  wire [15:0] _T_29198; // @[Mux.scala 19:72:@25318.4]
  wire [15:0] _T_29200; // @[Mux.scala 19:72:@25319.4]
  wire [7:0] _T_29207; // @[Mux.scala 19:72:@25326.4]
  wire [7:0] _T_29214; // @[Mux.scala 19:72:@25333.4]
  wire [15:0] _T_29215; // @[Mux.scala 19:72:@25334.4]
  wire [15:0] _T_29217; // @[Mux.scala 19:72:@25335.4]
  wire [7:0] _T_29224; // @[Mux.scala 19:72:@25342.4]
  wire [7:0] _T_29231; // @[Mux.scala 19:72:@25349.4]
  wire [15:0] _T_29232; // @[Mux.scala 19:72:@25350.4]
  wire [15:0] _T_29234; // @[Mux.scala 19:72:@25351.4]
  wire [7:0] _T_29241; // @[Mux.scala 19:72:@25358.4]
  wire [7:0] _T_29248; // @[Mux.scala 19:72:@25365.4]
  wire [15:0] _T_29249; // @[Mux.scala 19:72:@25366.4]
  wire [15:0] _T_29251; // @[Mux.scala 19:72:@25367.4]
  wire [7:0] _T_29258; // @[Mux.scala 19:72:@25374.4]
  wire [7:0] _T_29265; // @[Mux.scala 19:72:@25381.4]
  wire [15:0] _T_29266; // @[Mux.scala 19:72:@25382.4]
  wire [15:0] _T_29268; // @[Mux.scala 19:72:@25383.4]
  wire [7:0] _T_29275; // @[Mux.scala 19:72:@25390.4]
  wire [7:0] _T_29282; // @[Mux.scala 19:72:@25397.4]
  wire [15:0] _T_29283; // @[Mux.scala 19:72:@25398.4]
  wire [15:0] _T_29285; // @[Mux.scala 19:72:@25399.4]
  wire [15:0] _T_29300; // @[Mux.scala 19:72:@25414.4]
  wire [15:0] _T_29302; // @[Mux.scala 19:72:@25415.4]
  wire [15:0] _T_29317; // @[Mux.scala 19:72:@25430.4]
  wire [15:0] _T_29319; // @[Mux.scala 19:72:@25431.4]
  wire [15:0] _T_29334; // @[Mux.scala 19:72:@25446.4]
  wire [15:0] _T_29336; // @[Mux.scala 19:72:@25447.4]
  wire [15:0] _T_29351; // @[Mux.scala 19:72:@25462.4]
  wire [15:0] _T_29353; // @[Mux.scala 19:72:@25463.4]
  wire [15:0] _T_29368; // @[Mux.scala 19:72:@25478.4]
  wire [15:0] _T_29370; // @[Mux.scala 19:72:@25479.4]
  wire [15:0] _T_29385; // @[Mux.scala 19:72:@25494.4]
  wire [15:0] _T_29387; // @[Mux.scala 19:72:@25495.4]
  wire [15:0] _T_29402; // @[Mux.scala 19:72:@25510.4]
  wire [15:0] _T_29404; // @[Mux.scala 19:72:@25511.4]
  wire [15:0] _T_29419; // @[Mux.scala 19:72:@25526.4]
  wire [15:0] _T_29421; // @[Mux.scala 19:72:@25527.4]
  wire [15:0] _T_29422; // @[Mux.scala 19:72:@25528.4]
  wire [15:0] _T_29423; // @[Mux.scala 19:72:@25529.4]
  wire [15:0] _T_29424; // @[Mux.scala 19:72:@25530.4]
  wire [15:0] _T_29425; // @[Mux.scala 19:72:@25531.4]
  wire [15:0] _T_29426; // @[Mux.scala 19:72:@25532.4]
  wire [15:0] _T_29427; // @[Mux.scala 19:72:@25533.4]
  wire [15:0] _T_29428; // @[Mux.scala 19:72:@25534.4]
  wire [15:0] _T_29429; // @[Mux.scala 19:72:@25535.4]
  wire [15:0] _T_29430; // @[Mux.scala 19:72:@25536.4]
  wire [15:0] _T_29431; // @[Mux.scala 19:72:@25537.4]
  wire [15:0] _T_29432; // @[Mux.scala 19:72:@25538.4]
  wire [15:0] _T_29433; // @[Mux.scala 19:72:@25539.4]
  wire [15:0] _T_29434; // @[Mux.scala 19:72:@25540.4]
  wire [15:0] _T_29435; // @[Mux.scala 19:72:@25541.4]
  wire [15:0] _T_29436; // @[Mux.scala 19:72:@25542.4]
  wire [7:0] _T_30014; // @[Mux.scala 19:72:@25892.4]
  wire [7:0] _T_30021; // @[Mux.scala 19:72:@25899.4]
  wire [15:0] _T_30022; // @[Mux.scala 19:72:@25900.4]
  wire [15:0] _T_30024; // @[Mux.scala 19:72:@25901.4]
  wire [7:0] _T_30031; // @[Mux.scala 19:72:@25908.4]
  wire [7:0] _T_30038; // @[Mux.scala 19:72:@25915.4]
  wire [15:0] _T_30039; // @[Mux.scala 19:72:@25916.4]
  wire [15:0] _T_30041; // @[Mux.scala 19:72:@25917.4]
  wire [7:0] _T_30048; // @[Mux.scala 19:72:@25924.4]
  wire [7:0] _T_30055; // @[Mux.scala 19:72:@25931.4]
  wire [15:0] _T_30056; // @[Mux.scala 19:72:@25932.4]
  wire [15:0] _T_30058; // @[Mux.scala 19:72:@25933.4]
  wire [7:0] _T_30065; // @[Mux.scala 19:72:@25940.4]
  wire [7:0] _T_30072; // @[Mux.scala 19:72:@25947.4]
  wire [15:0] _T_30073; // @[Mux.scala 19:72:@25948.4]
  wire [15:0] _T_30075; // @[Mux.scala 19:72:@25949.4]
  wire [7:0] _T_30082; // @[Mux.scala 19:72:@25956.4]
  wire [7:0] _T_30089; // @[Mux.scala 19:72:@25963.4]
  wire [15:0] _T_30090; // @[Mux.scala 19:72:@25964.4]
  wire [15:0] _T_30092; // @[Mux.scala 19:72:@25965.4]
  wire [7:0] _T_30099; // @[Mux.scala 19:72:@25972.4]
  wire [7:0] _T_30106; // @[Mux.scala 19:72:@25979.4]
  wire [15:0] _T_30107; // @[Mux.scala 19:72:@25980.4]
  wire [15:0] _T_30109; // @[Mux.scala 19:72:@25981.4]
  wire [7:0] _T_30116; // @[Mux.scala 19:72:@25988.4]
  wire [7:0] _T_30123; // @[Mux.scala 19:72:@25995.4]
  wire [15:0] _T_30124; // @[Mux.scala 19:72:@25996.4]
  wire [15:0] _T_30126; // @[Mux.scala 19:72:@25997.4]
  wire [7:0] _T_30133; // @[Mux.scala 19:72:@26004.4]
  wire [7:0] _T_30140; // @[Mux.scala 19:72:@26011.4]
  wire [15:0] _T_30141; // @[Mux.scala 19:72:@26012.4]
  wire [15:0] _T_30143; // @[Mux.scala 19:72:@26013.4]
  wire [15:0] _T_30158; // @[Mux.scala 19:72:@26028.4]
  wire [15:0] _T_30160; // @[Mux.scala 19:72:@26029.4]
  wire [15:0] _T_30175; // @[Mux.scala 19:72:@26044.4]
  wire [15:0] _T_30177; // @[Mux.scala 19:72:@26045.4]
  wire [15:0] _T_30192; // @[Mux.scala 19:72:@26060.4]
  wire [15:0] _T_30194; // @[Mux.scala 19:72:@26061.4]
  wire [15:0] _T_30209; // @[Mux.scala 19:72:@26076.4]
  wire [15:0] _T_30211; // @[Mux.scala 19:72:@26077.4]
  wire [15:0] _T_30226; // @[Mux.scala 19:72:@26092.4]
  wire [15:0] _T_30228; // @[Mux.scala 19:72:@26093.4]
  wire [15:0] _T_30243; // @[Mux.scala 19:72:@26108.4]
  wire [15:0] _T_30245; // @[Mux.scala 19:72:@26109.4]
  wire [15:0] _T_30260; // @[Mux.scala 19:72:@26124.4]
  wire [15:0] _T_30262; // @[Mux.scala 19:72:@26125.4]
  wire [15:0] _T_30277; // @[Mux.scala 19:72:@26140.4]
  wire [15:0] _T_30279; // @[Mux.scala 19:72:@26141.4]
  wire [15:0] _T_30280; // @[Mux.scala 19:72:@26142.4]
  wire [15:0] _T_30281; // @[Mux.scala 19:72:@26143.4]
  wire [15:0] _T_30282; // @[Mux.scala 19:72:@26144.4]
  wire [15:0] _T_30283; // @[Mux.scala 19:72:@26145.4]
  wire [15:0] _T_30284; // @[Mux.scala 19:72:@26146.4]
  wire [15:0] _T_30285; // @[Mux.scala 19:72:@26147.4]
  wire [15:0] _T_30286; // @[Mux.scala 19:72:@26148.4]
  wire [15:0] _T_30287; // @[Mux.scala 19:72:@26149.4]
  wire [15:0] _T_30288; // @[Mux.scala 19:72:@26150.4]
  wire [15:0] _T_30289; // @[Mux.scala 19:72:@26151.4]
  wire [15:0] _T_30290; // @[Mux.scala 19:72:@26152.4]
  wire [15:0] _T_30291; // @[Mux.scala 19:72:@26153.4]
  wire [15:0] _T_30292; // @[Mux.scala 19:72:@26154.4]
  wire [15:0] _T_30293; // @[Mux.scala 19:72:@26155.4]
  wire [15:0] _T_30294; // @[Mux.scala 19:72:@26156.4]
  wire [7:0] _T_30872; // @[Mux.scala 19:72:@26506.4]
  wire [7:0] _T_30879; // @[Mux.scala 19:72:@26513.4]
  wire [15:0] _T_30880; // @[Mux.scala 19:72:@26514.4]
  wire [15:0] _T_30882; // @[Mux.scala 19:72:@26515.4]
  wire [7:0] _T_30889; // @[Mux.scala 19:72:@26522.4]
  wire [7:0] _T_30896; // @[Mux.scala 19:72:@26529.4]
  wire [15:0] _T_30897; // @[Mux.scala 19:72:@26530.4]
  wire [15:0] _T_30899; // @[Mux.scala 19:72:@26531.4]
  wire [7:0] _T_30906; // @[Mux.scala 19:72:@26538.4]
  wire [7:0] _T_30913; // @[Mux.scala 19:72:@26545.4]
  wire [15:0] _T_30914; // @[Mux.scala 19:72:@26546.4]
  wire [15:0] _T_30916; // @[Mux.scala 19:72:@26547.4]
  wire [7:0] _T_30923; // @[Mux.scala 19:72:@26554.4]
  wire [7:0] _T_30930; // @[Mux.scala 19:72:@26561.4]
  wire [15:0] _T_30931; // @[Mux.scala 19:72:@26562.4]
  wire [15:0] _T_30933; // @[Mux.scala 19:72:@26563.4]
  wire [7:0] _T_30940; // @[Mux.scala 19:72:@26570.4]
  wire [7:0] _T_30947; // @[Mux.scala 19:72:@26577.4]
  wire [15:0] _T_30948; // @[Mux.scala 19:72:@26578.4]
  wire [15:0] _T_30950; // @[Mux.scala 19:72:@26579.4]
  wire [7:0] _T_30957; // @[Mux.scala 19:72:@26586.4]
  wire [7:0] _T_30964; // @[Mux.scala 19:72:@26593.4]
  wire [15:0] _T_30965; // @[Mux.scala 19:72:@26594.4]
  wire [15:0] _T_30967; // @[Mux.scala 19:72:@26595.4]
  wire [7:0] _T_30974; // @[Mux.scala 19:72:@26602.4]
  wire [7:0] _T_30981; // @[Mux.scala 19:72:@26609.4]
  wire [15:0] _T_30982; // @[Mux.scala 19:72:@26610.4]
  wire [15:0] _T_30984; // @[Mux.scala 19:72:@26611.4]
  wire [7:0] _T_30991; // @[Mux.scala 19:72:@26618.4]
  wire [7:0] _T_30998; // @[Mux.scala 19:72:@26625.4]
  wire [15:0] _T_30999; // @[Mux.scala 19:72:@26626.4]
  wire [15:0] _T_31001; // @[Mux.scala 19:72:@26627.4]
  wire [15:0] _T_31016; // @[Mux.scala 19:72:@26642.4]
  wire [15:0] _T_31018; // @[Mux.scala 19:72:@26643.4]
  wire [15:0] _T_31033; // @[Mux.scala 19:72:@26658.4]
  wire [15:0] _T_31035; // @[Mux.scala 19:72:@26659.4]
  wire [15:0] _T_31050; // @[Mux.scala 19:72:@26674.4]
  wire [15:0] _T_31052; // @[Mux.scala 19:72:@26675.4]
  wire [15:0] _T_31067; // @[Mux.scala 19:72:@26690.4]
  wire [15:0] _T_31069; // @[Mux.scala 19:72:@26691.4]
  wire [15:0] _T_31084; // @[Mux.scala 19:72:@26706.4]
  wire [15:0] _T_31086; // @[Mux.scala 19:72:@26707.4]
  wire [15:0] _T_31101; // @[Mux.scala 19:72:@26722.4]
  wire [15:0] _T_31103; // @[Mux.scala 19:72:@26723.4]
  wire [15:0] _T_31118; // @[Mux.scala 19:72:@26738.4]
  wire [15:0] _T_31120; // @[Mux.scala 19:72:@26739.4]
  wire [15:0] _T_31135; // @[Mux.scala 19:72:@26754.4]
  wire [15:0] _T_31137; // @[Mux.scala 19:72:@26755.4]
  wire [15:0] _T_31138; // @[Mux.scala 19:72:@26756.4]
  wire [15:0] _T_31139; // @[Mux.scala 19:72:@26757.4]
  wire [15:0] _T_31140; // @[Mux.scala 19:72:@26758.4]
  wire [15:0] _T_31141; // @[Mux.scala 19:72:@26759.4]
  wire [15:0] _T_31142; // @[Mux.scala 19:72:@26760.4]
  wire [15:0] _T_31143; // @[Mux.scala 19:72:@26761.4]
  wire [15:0] _T_31144; // @[Mux.scala 19:72:@26762.4]
  wire [15:0] _T_31145; // @[Mux.scala 19:72:@26763.4]
  wire [15:0] _T_31146; // @[Mux.scala 19:72:@26764.4]
  wire [15:0] _T_31147; // @[Mux.scala 19:72:@26765.4]
  wire [15:0] _T_31148; // @[Mux.scala 19:72:@26766.4]
  wire [15:0] _T_31149; // @[Mux.scala 19:72:@26767.4]
  wire [15:0] _T_31150; // @[Mux.scala 19:72:@26768.4]
  wire [15:0] _T_31151; // @[Mux.scala 19:72:@26769.4]
  wire [15:0] _T_31152; // @[Mux.scala 19:72:@26770.4]
  reg  conflictPReg_0_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_163;
  reg  conflictPReg_0_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_164;
  reg  conflictPReg_0_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_165;
  reg  conflictPReg_0_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_166;
  reg  conflictPReg_0_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_167;
  reg  conflictPReg_0_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_168;
  reg  conflictPReg_0_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_169;
  reg  conflictPReg_0_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_170;
  reg  conflictPReg_0_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_171;
  reg  conflictPReg_0_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_172;
  reg  conflictPReg_0_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_173;
  reg  conflictPReg_0_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_174;
  reg  conflictPReg_0_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_175;
  reg  conflictPReg_0_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_176;
  reg  conflictPReg_0_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_177;
  reg  conflictPReg_0_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_178;
  reg  conflictPReg_1_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_179;
  reg  conflictPReg_1_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_180;
  reg  conflictPReg_1_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_181;
  reg  conflictPReg_1_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_182;
  reg  conflictPReg_1_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_183;
  reg  conflictPReg_1_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_184;
  reg  conflictPReg_1_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_185;
  reg  conflictPReg_1_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_186;
  reg  conflictPReg_1_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_187;
  reg  conflictPReg_1_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_188;
  reg  conflictPReg_1_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_189;
  reg  conflictPReg_1_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_190;
  reg  conflictPReg_1_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_191;
  reg  conflictPReg_1_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_192;
  reg  conflictPReg_1_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_193;
  reg  conflictPReg_1_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_194;
  reg  conflictPReg_2_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_195;
  reg  conflictPReg_2_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_196;
  reg  conflictPReg_2_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_197;
  reg  conflictPReg_2_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_198;
  reg  conflictPReg_2_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_199;
  reg  conflictPReg_2_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_200;
  reg  conflictPReg_2_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_201;
  reg  conflictPReg_2_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_202;
  reg  conflictPReg_2_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_203;
  reg  conflictPReg_2_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_204;
  reg  conflictPReg_2_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_205;
  reg  conflictPReg_2_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_206;
  reg  conflictPReg_2_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_207;
  reg  conflictPReg_2_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_208;
  reg  conflictPReg_2_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_209;
  reg  conflictPReg_2_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_210;
  reg  conflictPReg_3_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_211;
  reg  conflictPReg_3_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_212;
  reg  conflictPReg_3_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_213;
  reg  conflictPReg_3_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_214;
  reg  conflictPReg_3_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_215;
  reg  conflictPReg_3_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_216;
  reg  conflictPReg_3_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_217;
  reg  conflictPReg_3_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_218;
  reg  conflictPReg_3_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_219;
  reg  conflictPReg_3_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_220;
  reg  conflictPReg_3_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_221;
  reg  conflictPReg_3_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_222;
  reg  conflictPReg_3_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_223;
  reg  conflictPReg_3_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_224;
  reg  conflictPReg_3_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_225;
  reg  conflictPReg_3_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_226;
  reg  conflictPReg_4_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_227;
  reg  conflictPReg_4_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_228;
  reg  conflictPReg_4_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_229;
  reg  conflictPReg_4_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_230;
  reg  conflictPReg_4_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_231;
  reg  conflictPReg_4_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_232;
  reg  conflictPReg_4_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_233;
  reg  conflictPReg_4_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_234;
  reg  conflictPReg_4_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_235;
  reg  conflictPReg_4_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_236;
  reg  conflictPReg_4_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_237;
  reg  conflictPReg_4_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_238;
  reg  conflictPReg_4_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_239;
  reg  conflictPReg_4_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_240;
  reg  conflictPReg_4_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_241;
  reg  conflictPReg_4_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_242;
  reg  conflictPReg_5_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_243;
  reg  conflictPReg_5_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_244;
  reg  conflictPReg_5_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_245;
  reg  conflictPReg_5_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_246;
  reg  conflictPReg_5_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_247;
  reg  conflictPReg_5_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_248;
  reg  conflictPReg_5_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_249;
  reg  conflictPReg_5_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_250;
  reg  conflictPReg_5_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_251;
  reg  conflictPReg_5_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_252;
  reg  conflictPReg_5_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_253;
  reg  conflictPReg_5_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_254;
  reg  conflictPReg_5_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_255;
  reg  conflictPReg_5_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_256;
  reg  conflictPReg_5_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_257;
  reg  conflictPReg_5_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_258;
  reg  conflictPReg_6_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_259;
  reg  conflictPReg_6_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_260;
  reg  conflictPReg_6_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_261;
  reg  conflictPReg_6_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_262;
  reg  conflictPReg_6_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_263;
  reg  conflictPReg_6_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_264;
  reg  conflictPReg_6_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_265;
  reg  conflictPReg_6_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_266;
  reg  conflictPReg_6_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_267;
  reg  conflictPReg_6_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_268;
  reg  conflictPReg_6_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_269;
  reg  conflictPReg_6_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_270;
  reg  conflictPReg_6_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_271;
  reg  conflictPReg_6_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_272;
  reg  conflictPReg_6_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_273;
  reg  conflictPReg_6_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_274;
  reg  conflictPReg_7_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_275;
  reg  conflictPReg_7_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_276;
  reg  conflictPReg_7_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_277;
  reg  conflictPReg_7_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_278;
  reg  conflictPReg_7_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_279;
  reg  conflictPReg_7_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_280;
  reg  conflictPReg_7_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_281;
  reg  conflictPReg_7_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_282;
  reg  conflictPReg_7_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_283;
  reg  conflictPReg_7_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_284;
  reg  conflictPReg_7_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_285;
  reg  conflictPReg_7_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_286;
  reg  conflictPReg_7_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_287;
  reg  conflictPReg_7_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_288;
  reg  conflictPReg_7_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_289;
  reg  conflictPReg_7_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_290;
  reg  conflictPReg_8_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_291;
  reg  conflictPReg_8_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_292;
  reg  conflictPReg_8_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_293;
  reg  conflictPReg_8_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_294;
  reg  conflictPReg_8_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_295;
  reg  conflictPReg_8_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_296;
  reg  conflictPReg_8_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_297;
  reg  conflictPReg_8_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_298;
  reg  conflictPReg_8_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_299;
  reg  conflictPReg_8_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_300;
  reg  conflictPReg_8_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_301;
  reg  conflictPReg_8_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_302;
  reg  conflictPReg_8_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_303;
  reg  conflictPReg_8_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_304;
  reg  conflictPReg_8_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_305;
  reg  conflictPReg_8_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_306;
  reg  conflictPReg_9_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_307;
  reg  conflictPReg_9_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_308;
  reg  conflictPReg_9_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_309;
  reg  conflictPReg_9_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_310;
  reg  conflictPReg_9_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_311;
  reg  conflictPReg_9_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_312;
  reg  conflictPReg_9_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_313;
  reg  conflictPReg_9_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_314;
  reg  conflictPReg_9_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_315;
  reg  conflictPReg_9_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_316;
  reg  conflictPReg_9_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_317;
  reg  conflictPReg_9_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_318;
  reg  conflictPReg_9_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_319;
  reg  conflictPReg_9_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_320;
  reg  conflictPReg_9_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_321;
  reg  conflictPReg_9_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_322;
  reg  conflictPReg_10_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_323;
  reg  conflictPReg_10_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_324;
  reg  conflictPReg_10_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_325;
  reg  conflictPReg_10_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_326;
  reg  conflictPReg_10_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_327;
  reg  conflictPReg_10_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_328;
  reg  conflictPReg_10_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_329;
  reg  conflictPReg_10_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_330;
  reg  conflictPReg_10_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_331;
  reg  conflictPReg_10_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_332;
  reg  conflictPReg_10_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_333;
  reg  conflictPReg_10_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_334;
  reg  conflictPReg_10_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_335;
  reg  conflictPReg_10_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_336;
  reg  conflictPReg_10_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_337;
  reg  conflictPReg_10_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_338;
  reg  conflictPReg_11_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_339;
  reg  conflictPReg_11_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_340;
  reg  conflictPReg_11_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_341;
  reg  conflictPReg_11_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_342;
  reg  conflictPReg_11_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_343;
  reg  conflictPReg_11_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_344;
  reg  conflictPReg_11_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_345;
  reg  conflictPReg_11_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_346;
  reg  conflictPReg_11_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_347;
  reg  conflictPReg_11_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_348;
  reg  conflictPReg_11_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_349;
  reg  conflictPReg_11_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_350;
  reg  conflictPReg_11_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_351;
  reg  conflictPReg_11_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_352;
  reg  conflictPReg_11_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_353;
  reg  conflictPReg_11_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_354;
  reg  conflictPReg_12_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_355;
  reg  conflictPReg_12_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_356;
  reg  conflictPReg_12_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_357;
  reg  conflictPReg_12_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_358;
  reg  conflictPReg_12_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_359;
  reg  conflictPReg_12_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_360;
  reg  conflictPReg_12_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_361;
  reg  conflictPReg_12_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_362;
  reg  conflictPReg_12_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_363;
  reg  conflictPReg_12_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_364;
  reg  conflictPReg_12_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_365;
  reg  conflictPReg_12_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_366;
  reg  conflictPReg_12_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_367;
  reg  conflictPReg_12_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_368;
  reg  conflictPReg_12_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_369;
  reg  conflictPReg_12_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_370;
  reg  conflictPReg_13_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_371;
  reg  conflictPReg_13_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_372;
  reg  conflictPReg_13_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_373;
  reg  conflictPReg_13_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_374;
  reg  conflictPReg_13_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_375;
  reg  conflictPReg_13_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_376;
  reg  conflictPReg_13_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_377;
  reg  conflictPReg_13_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_378;
  reg  conflictPReg_13_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_379;
  reg  conflictPReg_13_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_380;
  reg  conflictPReg_13_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_381;
  reg  conflictPReg_13_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_382;
  reg  conflictPReg_13_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_383;
  reg  conflictPReg_13_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_384;
  reg  conflictPReg_13_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_385;
  reg  conflictPReg_13_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_386;
  reg  conflictPReg_14_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_387;
  reg  conflictPReg_14_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_388;
  reg  conflictPReg_14_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_389;
  reg  conflictPReg_14_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_390;
  reg  conflictPReg_14_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_391;
  reg  conflictPReg_14_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_392;
  reg  conflictPReg_14_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_393;
  reg  conflictPReg_14_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_394;
  reg  conflictPReg_14_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_395;
  reg  conflictPReg_14_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_396;
  reg  conflictPReg_14_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_397;
  reg  conflictPReg_14_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_398;
  reg  conflictPReg_14_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_399;
  reg  conflictPReg_14_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_400;
  reg  conflictPReg_14_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_401;
  reg  conflictPReg_14_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_402;
  reg  conflictPReg_15_0; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_403;
  reg  conflictPReg_15_1; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_404;
  reg  conflictPReg_15_2; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_405;
  reg  conflictPReg_15_3; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_406;
  reg  conflictPReg_15_4; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_407;
  reg  conflictPReg_15_5; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_408;
  reg  conflictPReg_15_6; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_409;
  reg  conflictPReg_15_7; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_410;
  reg  conflictPReg_15_8; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_411;
  reg  conflictPReg_15_9; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_412;
  reg  conflictPReg_15_10; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_413;
  reg  conflictPReg_15_11; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_414;
  reg  conflictPReg_15_12; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_415;
  reg  conflictPReg_15_13; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_416;
  reg  conflictPReg_15_14; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_417;
  reg  conflictPReg_15_15; // @[LoadQueue.scala 166:29:@27063.4]
  reg [31:0] _RAND_418;
  wire [7:0] _T_52326; // @[Mux.scala 19:72:@27634.4]
  wire [7:0] _T_52333; // @[Mux.scala 19:72:@27641.4]
  wire [15:0] _T_52334; // @[Mux.scala 19:72:@27642.4]
  wire [15:0] _T_52336; // @[Mux.scala 19:72:@27643.4]
  wire [7:0] _T_52343; // @[Mux.scala 19:72:@27650.4]
  wire [7:0] _T_52350; // @[Mux.scala 19:72:@27657.4]
  wire [15:0] _T_52351; // @[Mux.scala 19:72:@27658.4]
  wire [15:0] _T_52353; // @[Mux.scala 19:72:@27659.4]
  wire [7:0] _T_52360; // @[Mux.scala 19:72:@27666.4]
  wire [7:0] _T_52367; // @[Mux.scala 19:72:@27673.4]
  wire [15:0] _T_52368; // @[Mux.scala 19:72:@27674.4]
  wire [15:0] _T_52370; // @[Mux.scala 19:72:@27675.4]
  wire [7:0] _T_52377; // @[Mux.scala 19:72:@27682.4]
  wire [7:0] _T_52384; // @[Mux.scala 19:72:@27689.4]
  wire [15:0] _T_52385; // @[Mux.scala 19:72:@27690.4]
  wire [15:0] _T_52387; // @[Mux.scala 19:72:@27691.4]
  wire [7:0] _T_52394; // @[Mux.scala 19:72:@27698.4]
  wire [7:0] _T_52401; // @[Mux.scala 19:72:@27705.4]
  wire [15:0] _T_52402; // @[Mux.scala 19:72:@27706.4]
  wire [15:0] _T_52404; // @[Mux.scala 19:72:@27707.4]
  wire [7:0] _T_52411; // @[Mux.scala 19:72:@27714.4]
  wire [7:0] _T_52418; // @[Mux.scala 19:72:@27721.4]
  wire [15:0] _T_52419; // @[Mux.scala 19:72:@27722.4]
  wire [15:0] _T_52421; // @[Mux.scala 19:72:@27723.4]
  wire [7:0] _T_52428; // @[Mux.scala 19:72:@27730.4]
  wire [7:0] _T_52435; // @[Mux.scala 19:72:@27737.4]
  wire [15:0] _T_52436; // @[Mux.scala 19:72:@27738.4]
  wire [15:0] _T_52438; // @[Mux.scala 19:72:@27739.4]
  wire [7:0] _T_52445; // @[Mux.scala 19:72:@27746.4]
  wire [7:0] _T_52452; // @[Mux.scala 19:72:@27753.4]
  wire [15:0] _T_52453; // @[Mux.scala 19:72:@27754.4]
  wire [15:0] _T_52455; // @[Mux.scala 19:72:@27755.4]
  wire [15:0] _T_52470; // @[Mux.scala 19:72:@27770.4]
  wire [15:0] _T_52472; // @[Mux.scala 19:72:@27771.4]
  wire [15:0] _T_52487; // @[Mux.scala 19:72:@27786.4]
  wire [15:0] _T_52489; // @[Mux.scala 19:72:@27787.4]
  wire [15:0] _T_52504; // @[Mux.scala 19:72:@27802.4]
  wire [15:0] _T_52506; // @[Mux.scala 19:72:@27803.4]
  wire [15:0] _T_52521; // @[Mux.scala 19:72:@27818.4]
  wire [15:0] _T_52523; // @[Mux.scala 19:72:@27819.4]
  wire [15:0] _T_52538; // @[Mux.scala 19:72:@27834.4]
  wire [15:0] _T_52540; // @[Mux.scala 19:72:@27835.4]
  wire [15:0] _T_52555; // @[Mux.scala 19:72:@27850.4]
  wire [15:0] _T_52557; // @[Mux.scala 19:72:@27851.4]
  wire [15:0] _T_52572; // @[Mux.scala 19:72:@27866.4]
  wire [15:0] _T_52574; // @[Mux.scala 19:72:@27867.4]
  wire [15:0] _T_52589; // @[Mux.scala 19:72:@27882.4]
  wire [15:0] _T_52591; // @[Mux.scala 19:72:@27883.4]
  wire [15:0] _T_52592; // @[Mux.scala 19:72:@27884.4]
  wire [15:0] _T_52593; // @[Mux.scala 19:72:@27885.4]
  wire [15:0] _T_52594; // @[Mux.scala 19:72:@27886.4]
  wire [15:0] _T_52595; // @[Mux.scala 19:72:@27887.4]
  wire [15:0] _T_52596; // @[Mux.scala 19:72:@27888.4]
  wire [15:0] _T_52597; // @[Mux.scala 19:72:@27889.4]
  wire [15:0] _T_52598; // @[Mux.scala 19:72:@27890.4]
  wire [15:0] _T_52599; // @[Mux.scala 19:72:@27891.4]
  wire [15:0] _T_52600; // @[Mux.scala 19:72:@27892.4]
  wire [15:0] _T_52601; // @[Mux.scala 19:72:@27893.4]
  wire [15:0] _T_52602; // @[Mux.scala 19:72:@27894.4]
  wire [15:0] _T_52603; // @[Mux.scala 19:72:@27895.4]
  wire [15:0] _T_52604; // @[Mux.scala 19:72:@27896.4]
  wire [15:0] _T_52605; // @[Mux.scala 19:72:@27897.4]
  wire [15:0] _T_52606; // @[Mux.scala 19:72:@27898.4]
  wire [7:0] _T_53184; // @[Mux.scala 19:72:@28248.4]
  wire [7:0] _T_53191; // @[Mux.scala 19:72:@28255.4]
  wire [15:0] _T_53192; // @[Mux.scala 19:72:@28256.4]
  wire [15:0] _T_53194; // @[Mux.scala 19:72:@28257.4]
  wire [7:0] _T_53201; // @[Mux.scala 19:72:@28264.4]
  wire [7:0] _T_53208; // @[Mux.scala 19:72:@28271.4]
  wire [15:0] _T_53209; // @[Mux.scala 19:72:@28272.4]
  wire [15:0] _T_53211; // @[Mux.scala 19:72:@28273.4]
  wire [7:0] _T_53218; // @[Mux.scala 19:72:@28280.4]
  wire [7:0] _T_53225; // @[Mux.scala 19:72:@28287.4]
  wire [15:0] _T_53226; // @[Mux.scala 19:72:@28288.4]
  wire [15:0] _T_53228; // @[Mux.scala 19:72:@28289.4]
  wire [7:0] _T_53235; // @[Mux.scala 19:72:@28296.4]
  wire [7:0] _T_53242; // @[Mux.scala 19:72:@28303.4]
  wire [15:0] _T_53243; // @[Mux.scala 19:72:@28304.4]
  wire [15:0] _T_53245; // @[Mux.scala 19:72:@28305.4]
  wire [7:0] _T_53252; // @[Mux.scala 19:72:@28312.4]
  wire [7:0] _T_53259; // @[Mux.scala 19:72:@28319.4]
  wire [15:0] _T_53260; // @[Mux.scala 19:72:@28320.4]
  wire [15:0] _T_53262; // @[Mux.scala 19:72:@28321.4]
  wire [7:0] _T_53269; // @[Mux.scala 19:72:@28328.4]
  wire [7:0] _T_53276; // @[Mux.scala 19:72:@28335.4]
  wire [15:0] _T_53277; // @[Mux.scala 19:72:@28336.4]
  wire [15:0] _T_53279; // @[Mux.scala 19:72:@28337.4]
  wire [7:0] _T_53286; // @[Mux.scala 19:72:@28344.4]
  wire [7:0] _T_53293; // @[Mux.scala 19:72:@28351.4]
  wire [15:0] _T_53294; // @[Mux.scala 19:72:@28352.4]
  wire [15:0] _T_53296; // @[Mux.scala 19:72:@28353.4]
  wire [7:0] _T_53303; // @[Mux.scala 19:72:@28360.4]
  wire [7:0] _T_53310; // @[Mux.scala 19:72:@28367.4]
  wire [15:0] _T_53311; // @[Mux.scala 19:72:@28368.4]
  wire [15:0] _T_53313; // @[Mux.scala 19:72:@28369.4]
  wire [15:0] _T_53328; // @[Mux.scala 19:72:@28384.4]
  wire [15:0] _T_53330; // @[Mux.scala 19:72:@28385.4]
  wire [15:0] _T_53345; // @[Mux.scala 19:72:@28400.4]
  wire [15:0] _T_53347; // @[Mux.scala 19:72:@28401.4]
  wire [15:0] _T_53362; // @[Mux.scala 19:72:@28416.4]
  wire [15:0] _T_53364; // @[Mux.scala 19:72:@28417.4]
  wire [15:0] _T_53379; // @[Mux.scala 19:72:@28432.4]
  wire [15:0] _T_53381; // @[Mux.scala 19:72:@28433.4]
  wire [15:0] _T_53396; // @[Mux.scala 19:72:@28448.4]
  wire [15:0] _T_53398; // @[Mux.scala 19:72:@28449.4]
  wire [15:0] _T_53413; // @[Mux.scala 19:72:@28464.4]
  wire [15:0] _T_53415; // @[Mux.scala 19:72:@28465.4]
  wire [15:0] _T_53430; // @[Mux.scala 19:72:@28480.4]
  wire [15:0] _T_53432; // @[Mux.scala 19:72:@28481.4]
  wire [15:0] _T_53447; // @[Mux.scala 19:72:@28496.4]
  wire [15:0] _T_53449; // @[Mux.scala 19:72:@28497.4]
  wire [15:0] _T_53450; // @[Mux.scala 19:72:@28498.4]
  wire [15:0] _T_53451; // @[Mux.scala 19:72:@28499.4]
  wire [15:0] _T_53452; // @[Mux.scala 19:72:@28500.4]
  wire [15:0] _T_53453; // @[Mux.scala 19:72:@28501.4]
  wire [15:0] _T_53454; // @[Mux.scala 19:72:@28502.4]
  wire [15:0] _T_53455; // @[Mux.scala 19:72:@28503.4]
  wire [15:0] _T_53456; // @[Mux.scala 19:72:@28504.4]
  wire [15:0] _T_53457; // @[Mux.scala 19:72:@28505.4]
  wire [15:0] _T_53458; // @[Mux.scala 19:72:@28506.4]
  wire [15:0] _T_53459; // @[Mux.scala 19:72:@28507.4]
  wire [15:0] _T_53460; // @[Mux.scala 19:72:@28508.4]
  wire [15:0] _T_53461; // @[Mux.scala 19:72:@28509.4]
  wire [15:0] _T_53462; // @[Mux.scala 19:72:@28510.4]
  wire [15:0] _T_53463; // @[Mux.scala 19:72:@28511.4]
  wire [15:0] _T_53464; // @[Mux.scala 19:72:@28512.4]
  wire [7:0] _T_54042; // @[Mux.scala 19:72:@28862.4]
  wire [7:0] _T_54049; // @[Mux.scala 19:72:@28869.4]
  wire [15:0] _T_54050; // @[Mux.scala 19:72:@28870.4]
  wire [15:0] _T_54052; // @[Mux.scala 19:72:@28871.4]
  wire [7:0] _T_54059; // @[Mux.scala 19:72:@28878.4]
  wire [7:0] _T_54066; // @[Mux.scala 19:72:@28885.4]
  wire [15:0] _T_54067; // @[Mux.scala 19:72:@28886.4]
  wire [15:0] _T_54069; // @[Mux.scala 19:72:@28887.4]
  wire [7:0] _T_54076; // @[Mux.scala 19:72:@28894.4]
  wire [7:0] _T_54083; // @[Mux.scala 19:72:@28901.4]
  wire [15:0] _T_54084; // @[Mux.scala 19:72:@28902.4]
  wire [15:0] _T_54086; // @[Mux.scala 19:72:@28903.4]
  wire [7:0] _T_54093; // @[Mux.scala 19:72:@28910.4]
  wire [7:0] _T_54100; // @[Mux.scala 19:72:@28917.4]
  wire [15:0] _T_54101; // @[Mux.scala 19:72:@28918.4]
  wire [15:0] _T_54103; // @[Mux.scala 19:72:@28919.4]
  wire [7:0] _T_54110; // @[Mux.scala 19:72:@28926.4]
  wire [7:0] _T_54117; // @[Mux.scala 19:72:@28933.4]
  wire [15:0] _T_54118; // @[Mux.scala 19:72:@28934.4]
  wire [15:0] _T_54120; // @[Mux.scala 19:72:@28935.4]
  wire [7:0] _T_54127; // @[Mux.scala 19:72:@28942.4]
  wire [7:0] _T_54134; // @[Mux.scala 19:72:@28949.4]
  wire [15:0] _T_54135; // @[Mux.scala 19:72:@28950.4]
  wire [15:0] _T_54137; // @[Mux.scala 19:72:@28951.4]
  wire [7:0] _T_54144; // @[Mux.scala 19:72:@28958.4]
  wire [7:0] _T_54151; // @[Mux.scala 19:72:@28965.4]
  wire [15:0] _T_54152; // @[Mux.scala 19:72:@28966.4]
  wire [15:0] _T_54154; // @[Mux.scala 19:72:@28967.4]
  wire [7:0] _T_54161; // @[Mux.scala 19:72:@28974.4]
  wire [7:0] _T_54168; // @[Mux.scala 19:72:@28981.4]
  wire [15:0] _T_54169; // @[Mux.scala 19:72:@28982.4]
  wire [15:0] _T_54171; // @[Mux.scala 19:72:@28983.4]
  wire [15:0] _T_54186; // @[Mux.scala 19:72:@28998.4]
  wire [15:0] _T_54188; // @[Mux.scala 19:72:@28999.4]
  wire [15:0] _T_54203; // @[Mux.scala 19:72:@29014.4]
  wire [15:0] _T_54205; // @[Mux.scala 19:72:@29015.4]
  wire [15:0] _T_54220; // @[Mux.scala 19:72:@29030.4]
  wire [15:0] _T_54222; // @[Mux.scala 19:72:@29031.4]
  wire [15:0] _T_54237; // @[Mux.scala 19:72:@29046.4]
  wire [15:0] _T_54239; // @[Mux.scala 19:72:@29047.4]
  wire [15:0] _T_54254; // @[Mux.scala 19:72:@29062.4]
  wire [15:0] _T_54256; // @[Mux.scala 19:72:@29063.4]
  wire [15:0] _T_54271; // @[Mux.scala 19:72:@29078.4]
  wire [15:0] _T_54273; // @[Mux.scala 19:72:@29079.4]
  wire [15:0] _T_54288; // @[Mux.scala 19:72:@29094.4]
  wire [15:0] _T_54290; // @[Mux.scala 19:72:@29095.4]
  wire [15:0] _T_54305; // @[Mux.scala 19:72:@29110.4]
  wire [15:0] _T_54307; // @[Mux.scala 19:72:@29111.4]
  wire [15:0] _T_54308; // @[Mux.scala 19:72:@29112.4]
  wire [15:0] _T_54309; // @[Mux.scala 19:72:@29113.4]
  wire [15:0] _T_54310; // @[Mux.scala 19:72:@29114.4]
  wire [15:0] _T_54311; // @[Mux.scala 19:72:@29115.4]
  wire [15:0] _T_54312; // @[Mux.scala 19:72:@29116.4]
  wire [15:0] _T_54313; // @[Mux.scala 19:72:@29117.4]
  wire [15:0] _T_54314; // @[Mux.scala 19:72:@29118.4]
  wire [15:0] _T_54315; // @[Mux.scala 19:72:@29119.4]
  wire [15:0] _T_54316; // @[Mux.scala 19:72:@29120.4]
  wire [15:0] _T_54317; // @[Mux.scala 19:72:@29121.4]
  wire [15:0] _T_54318; // @[Mux.scala 19:72:@29122.4]
  wire [15:0] _T_54319; // @[Mux.scala 19:72:@29123.4]
  wire [15:0] _T_54320; // @[Mux.scala 19:72:@29124.4]
  wire [15:0] _T_54321; // @[Mux.scala 19:72:@29125.4]
  wire [15:0] _T_54322; // @[Mux.scala 19:72:@29126.4]
  wire [7:0] _T_54900; // @[Mux.scala 19:72:@29476.4]
  wire [7:0] _T_54907; // @[Mux.scala 19:72:@29483.4]
  wire [15:0] _T_54908; // @[Mux.scala 19:72:@29484.4]
  wire [15:0] _T_54910; // @[Mux.scala 19:72:@29485.4]
  wire [7:0] _T_54917; // @[Mux.scala 19:72:@29492.4]
  wire [7:0] _T_54924; // @[Mux.scala 19:72:@29499.4]
  wire [15:0] _T_54925; // @[Mux.scala 19:72:@29500.4]
  wire [15:0] _T_54927; // @[Mux.scala 19:72:@29501.4]
  wire [7:0] _T_54934; // @[Mux.scala 19:72:@29508.4]
  wire [7:0] _T_54941; // @[Mux.scala 19:72:@29515.4]
  wire [15:0] _T_54942; // @[Mux.scala 19:72:@29516.4]
  wire [15:0] _T_54944; // @[Mux.scala 19:72:@29517.4]
  wire [7:0] _T_54951; // @[Mux.scala 19:72:@29524.4]
  wire [7:0] _T_54958; // @[Mux.scala 19:72:@29531.4]
  wire [15:0] _T_54959; // @[Mux.scala 19:72:@29532.4]
  wire [15:0] _T_54961; // @[Mux.scala 19:72:@29533.4]
  wire [7:0] _T_54968; // @[Mux.scala 19:72:@29540.4]
  wire [7:0] _T_54975; // @[Mux.scala 19:72:@29547.4]
  wire [15:0] _T_54976; // @[Mux.scala 19:72:@29548.4]
  wire [15:0] _T_54978; // @[Mux.scala 19:72:@29549.4]
  wire [7:0] _T_54985; // @[Mux.scala 19:72:@29556.4]
  wire [7:0] _T_54992; // @[Mux.scala 19:72:@29563.4]
  wire [15:0] _T_54993; // @[Mux.scala 19:72:@29564.4]
  wire [15:0] _T_54995; // @[Mux.scala 19:72:@29565.4]
  wire [7:0] _T_55002; // @[Mux.scala 19:72:@29572.4]
  wire [7:0] _T_55009; // @[Mux.scala 19:72:@29579.4]
  wire [15:0] _T_55010; // @[Mux.scala 19:72:@29580.4]
  wire [15:0] _T_55012; // @[Mux.scala 19:72:@29581.4]
  wire [7:0] _T_55019; // @[Mux.scala 19:72:@29588.4]
  wire [7:0] _T_55026; // @[Mux.scala 19:72:@29595.4]
  wire [15:0] _T_55027; // @[Mux.scala 19:72:@29596.4]
  wire [15:0] _T_55029; // @[Mux.scala 19:72:@29597.4]
  wire [15:0] _T_55044; // @[Mux.scala 19:72:@29612.4]
  wire [15:0] _T_55046; // @[Mux.scala 19:72:@29613.4]
  wire [15:0] _T_55061; // @[Mux.scala 19:72:@29628.4]
  wire [15:0] _T_55063; // @[Mux.scala 19:72:@29629.4]
  wire [15:0] _T_55078; // @[Mux.scala 19:72:@29644.4]
  wire [15:0] _T_55080; // @[Mux.scala 19:72:@29645.4]
  wire [15:0] _T_55095; // @[Mux.scala 19:72:@29660.4]
  wire [15:0] _T_55097; // @[Mux.scala 19:72:@29661.4]
  wire [15:0] _T_55112; // @[Mux.scala 19:72:@29676.4]
  wire [15:0] _T_55114; // @[Mux.scala 19:72:@29677.4]
  wire [15:0] _T_55129; // @[Mux.scala 19:72:@29692.4]
  wire [15:0] _T_55131; // @[Mux.scala 19:72:@29693.4]
  wire [15:0] _T_55146; // @[Mux.scala 19:72:@29708.4]
  wire [15:0] _T_55148; // @[Mux.scala 19:72:@29709.4]
  wire [15:0] _T_55163; // @[Mux.scala 19:72:@29724.4]
  wire [15:0] _T_55165; // @[Mux.scala 19:72:@29725.4]
  wire [15:0] _T_55166; // @[Mux.scala 19:72:@29726.4]
  wire [15:0] _T_55167; // @[Mux.scala 19:72:@29727.4]
  wire [15:0] _T_55168; // @[Mux.scala 19:72:@29728.4]
  wire [15:0] _T_55169; // @[Mux.scala 19:72:@29729.4]
  wire [15:0] _T_55170; // @[Mux.scala 19:72:@29730.4]
  wire [15:0] _T_55171; // @[Mux.scala 19:72:@29731.4]
  wire [15:0] _T_55172; // @[Mux.scala 19:72:@29732.4]
  wire [15:0] _T_55173; // @[Mux.scala 19:72:@29733.4]
  wire [15:0] _T_55174; // @[Mux.scala 19:72:@29734.4]
  wire [15:0] _T_55175; // @[Mux.scala 19:72:@29735.4]
  wire [15:0] _T_55176; // @[Mux.scala 19:72:@29736.4]
  wire [15:0] _T_55177; // @[Mux.scala 19:72:@29737.4]
  wire [15:0] _T_55178; // @[Mux.scala 19:72:@29738.4]
  wire [15:0] _T_55179; // @[Mux.scala 19:72:@29739.4]
  wire [15:0] _T_55180; // @[Mux.scala 19:72:@29740.4]
  wire [7:0] _T_55758; // @[Mux.scala 19:72:@30090.4]
  wire [7:0] _T_55765; // @[Mux.scala 19:72:@30097.4]
  wire [15:0] _T_55766; // @[Mux.scala 19:72:@30098.4]
  wire [15:0] _T_55768; // @[Mux.scala 19:72:@30099.4]
  wire [7:0] _T_55775; // @[Mux.scala 19:72:@30106.4]
  wire [7:0] _T_55782; // @[Mux.scala 19:72:@30113.4]
  wire [15:0] _T_55783; // @[Mux.scala 19:72:@30114.4]
  wire [15:0] _T_55785; // @[Mux.scala 19:72:@30115.4]
  wire [7:0] _T_55792; // @[Mux.scala 19:72:@30122.4]
  wire [7:0] _T_55799; // @[Mux.scala 19:72:@30129.4]
  wire [15:0] _T_55800; // @[Mux.scala 19:72:@30130.4]
  wire [15:0] _T_55802; // @[Mux.scala 19:72:@30131.4]
  wire [7:0] _T_55809; // @[Mux.scala 19:72:@30138.4]
  wire [7:0] _T_55816; // @[Mux.scala 19:72:@30145.4]
  wire [15:0] _T_55817; // @[Mux.scala 19:72:@30146.4]
  wire [15:0] _T_55819; // @[Mux.scala 19:72:@30147.4]
  wire [7:0] _T_55826; // @[Mux.scala 19:72:@30154.4]
  wire [7:0] _T_55833; // @[Mux.scala 19:72:@30161.4]
  wire [15:0] _T_55834; // @[Mux.scala 19:72:@30162.4]
  wire [15:0] _T_55836; // @[Mux.scala 19:72:@30163.4]
  wire [7:0] _T_55843; // @[Mux.scala 19:72:@30170.4]
  wire [7:0] _T_55850; // @[Mux.scala 19:72:@30177.4]
  wire [15:0] _T_55851; // @[Mux.scala 19:72:@30178.4]
  wire [15:0] _T_55853; // @[Mux.scala 19:72:@30179.4]
  wire [7:0] _T_55860; // @[Mux.scala 19:72:@30186.4]
  wire [7:0] _T_55867; // @[Mux.scala 19:72:@30193.4]
  wire [15:0] _T_55868; // @[Mux.scala 19:72:@30194.4]
  wire [15:0] _T_55870; // @[Mux.scala 19:72:@30195.4]
  wire [7:0] _T_55877; // @[Mux.scala 19:72:@30202.4]
  wire [7:0] _T_55884; // @[Mux.scala 19:72:@30209.4]
  wire [15:0] _T_55885; // @[Mux.scala 19:72:@30210.4]
  wire [15:0] _T_55887; // @[Mux.scala 19:72:@30211.4]
  wire [15:0] _T_55902; // @[Mux.scala 19:72:@30226.4]
  wire [15:0] _T_55904; // @[Mux.scala 19:72:@30227.4]
  wire [15:0] _T_55919; // @[Mux.scala 19:72:@30242.4]
  wire [15:0] _T_55921; // @[Mux.scala 19:72:@30243.4]
  wire [15:0] _T_55936; // @[Mux.scala 19:72:@30258.4]
  wire [15:0] _T_55938; // @[Mux.scala 19:72:@30259.4]
  wire [15:0] _T_55953; // @[Mux.scala 19:72:@30274.4]
  wire [15:0] _T_55955; // @[Mux.scala 19:72:@30275.4]
  wire [15:0] _T_55970; // @[Mux.scala 19:72:@30290.4]
  wire [15:0] _T_55972; // @[Mux.scala 19:72:@30291.4]
  wire [15:0] _T_55987; // @[Mux.scala 19:72:@30306.4]
  wire [15:0] _T_55989; // @[Mux.scala 19:72:@30307.4]
  wire [15:0] _T_56004; // @[Mux.scala 19:72:@30322.4]
  wire [15:0] _T_56006; // @[Mux.scala 19:72:@30323.4]
  wire [15:0] _T_56021; // @[Mux.scala 19:72:@30338.4]
  wire [15:0] _T_56023; // @[Mux.scala 19:72:@30339.4]
  wire [15:0] _T_56024; // @[Mux.scala 19:72:@30340.4]
  wire [15:0] _T_56025; // @[Mux.scala 19:72:@30341.4]
  wire [15:0] _T_56026; // @[Mux.scala 19:72:@30342.4]
  wire [15:0] _T_56027; // @[Mux.scala 19:72:@30343.4]
  wire [15:0] _T_56028; // @[Mux.scala 19:72:@30344.4]
  wire [15:0] _T_56029; // @[Mux.scala 19:72:@30345.4]
  wire [15:0] _T_56030; // @[Mux.scala 19:72:@30346.4]
  wire [15:0] _T_56031; // @[Mux.scala 19:72:@30347.4]
  wire [15:0] _T_56032; // @[Mux.scala 19:72:@30348.4]
  wire [15:0] _T_56033; // @[Mux.scala 19:72:@30349.4]
  wire [15:0] _T_56034; // @[Mux.scala 19:72:@30350.4]
  wire [15:0] _T_56035; // @[Mux.scala 19:72:@30351.4]
  wire [15:0] _T_56036; // @[Mux.scala 19:72:@30352.4]
  wire [15:0] _T_56037; // @[Mux.scala 19:72:@30353.4]
  wire [15:0] _T_56038; // @[Mux.scala 19:72:@30354.4]
  wire [7:0] _T_56616; // @[Mux.scala 19:72:@30704.4]
  wire [7:0] _T_56623; // @[Mux.scala 19:72:@30711.4]
  wire [15:0] _T_56624; // @[Mux.scala 19:72:@30712.4]
  wire [15:0] _T_56626; // @[Mux.scala 19:72:@30713.4]
  wire [7:0] _T_56633; // @[Mux.scala 19:72:@30720.4]
  wire [7:0] _T_56640; // @[Mux.scala 19:72:@30727.4]
  wire [15:0] _T_56641; // @[Mux.scala 19:72:@30728.4]
  wire [15:0] _T_56643; // @[Mux.scala 19:72:@30729.4]
  wire [7:0] _T_56650; // @[Mux.scala 19:72:@30736.4]
  wire [7:0] _T_56657; // @[Mux.scala 19:72:@30743.4]
  wire [15:0] _T_56658; // @[Mux.scala 19:72:@30744.4]
  wire [15:0] _T_56660; // @[Mux.scala 19:72:@30745.4]
  wire [7:0] _T_56667; // @[Mux.scala 19:72:@30752.4]
  wire [7:0] _T_56674; // @[Mux.scala 19:72:@30759.4]
  wire [15:0] _T_56675; // @[Mux.scala 19:72:@30760.4]
  wire [15:0] _T_56677; // @[Mux.scala 19:72:@30761.4]
  wire [7:0] _T_56684; // @[Mux.scala 19:72:@30768.4]
  wire [7:0] _T_56691; // @[Mux.scala 19:72:@30775.4]
  wire [15:0] _T_56692; // @[Mux.scala 19:72:@30776.4]
  wire [15:0] _T_56694; // @[Mux.scala 19:72:@30777.4]
  wire [7:0] _T_56701; // @[Mux.scala 19:72:@30784.4]
  wire [7:0] _T_56708; // @[Mux.scala 19:72:@30791.4]
  wire [15:0] _T_56709; // @[Mux.scala 19:72:@30792.4]
  wire [15:0] _T_56711; // @[Mux.scala 19:72:@30793.4]
  wire [7:0] _T_56718; // @[Mux.scala 19:72:@30800.4]
  wire [7:0] _T_56725; // @[Mux.scala 19:72:@30807.4]
  wire [15:0] _T_56726; // @[Mux.scala 19:72:@30808.4]
  wire [15:0] _T_56728; // @[Mux.scala 19:72:@30809.4]
  wire [7:0] _T_56735; // @[Mux.scala 19:72:@30816.4]
  wire [7:0] _T_56742; // @[Mux.scala 19:72:@30823.4]
  wire [15:0] _T_56743; // @[Mux.scala 19:72:@30824.4]
  wire [15:0] _T_56745; // @[Mux.scala 19:72:@30825.4]
  wire [15:0] _T_56760; // @[Mux.scala 19:72:@30840.4]
  wire [15:0] _T_56762; // @[Mux.scala 19:72:@30841.4]
  wire [15:0] _T_56777; // @[Mux.scala 19:72:@30856.4]
  wire [15:0] _T_56779; // @[Mux.scala 19:72:@30857.4]
  wire [15:0] _T_56794; // @[Mux.scala 19:72:@30872.4]
  wire [15:0] _T_56796; // @[Mux.scala 19:72:@30873.4]
  wire [15:0] _T_56811; // @[Mux.scala 19:72:@30888.4]
  wire [15:0] _T_56813; // @[Mux.scala 19:72:@30889.4]
  wire [15:0] _T_56828; // @[Mux.scala 19:72:@30904.4]
  wire [15:0] _T_56830; // @[Mux.scala 19:72:@30905.4]
  wire [15:0] _T_56845; // @[Mux.scala 19:72:@30920.4]
  wire [15:0] _T_56847; // @[Mux.scala 19:72:@30921.4]
  wire [15:0] _T_56862; // @[Mux.scala 19:72:@30936.4]
  wire [15:0] _T_56864; // @[Mux.scala 19:72:@30937.4]
  wire [15:0] _T_56879; // @[Mux.scala 19:72:@30952.4]
  wire [15:0] _T_56881; // @[Mux.scala 19:72:@30953.4]
  wire [15:0] _T_56882; // @[Mux.scala 19:72:@30954.4]
  wire [15:0] _T_56883; // @[Mux.scala 19:72:@30955.4]
  wire [15:0] _T_56884; // @[Mux.scala 19:72:@30956.4]
  wire [15:0] _T_56885; // @[Mux.scala 19:72:@30957.4]
  wire [15:0] _T_56886; // @[Mux.scala 19:72:@30958.4]
  wire [15:0] _T_56887; // @[Mux.scala 19:72:@30959.4]
  wire [15:0] _T_56888; // @[Mux.scala 19:72:@30960.4]
  wire [15:0] _T_56889; // @[Mux.scala 19:72:@30961.4]
  wire [15:0] _T_56890; // @[Mux.scala 19:72:@30962.4]
  wire [15:0] _T_56891; // @[Mux.scala 19:72:@30963.4]
  wire [15:0] _T_56892; // @[Mux.scala 19:72:@30964.4]
  wire [15:0] _T_56893; // @[Mux.scala 19:72:@30965.4]
  wire [15:0] _T_56894; // @[Mux.scala 19:72:@30966.4]
  wire [15:0] _T_56895; // @[Mux.scala 19:72:@30967.4]
  wire [15:0] _T_56896; // @[Mux.scala 19:72:@30968.4]
  wire [7:0] _T_57474; // @[Mux.scala 19:72:@31318.4]
  wire [7:0] _T_57481; // @[Mux.scala 19:72:@31325.4]
  wire [15:0] _T_57482; // @[Mux.scala 19:72:@31326.4]
  wire [15:0] _T_57484; // @[Mux.scala 19:72:@31327.4]
  wire [7:0] _T_57491; // @[Mux.scala 19:72:@31334.4]
  wire [7:0] _T_57498; // @[Mux.scala 19:72:@31341.4]
  wire [15:0] _T_57499; // @[Mux.scala 19:72:@31342.4]
  wire [15:0] _T_57501; // @[Mux.scala 19:72:@31343.4]
  wire [7:0] _T_57508; // @[Mux.scala 19:72:@31350.4]
  wire [7:0] _T_57515; // @[Mux.scala 19:72:@31357.4]
  wire [15:0] _T_57516; // @[Mux.scala 19:72:@31358.4]
  wire [15:0] _T_57518; // @[Mux.scala 19:72:@31359.4]
  wire [7:0] _T_57525; // @[Mux.scala 19:72:@31366.4]
  wire [7:0] _T_57532; // @[Mux.scala 19:72:@31373.4]
  wire [15:0] _T_57533; // @[Mux.scala 19:72:@31374.4]
  wire [15:0] _T_57535; // @[Mux.scala 19:72:@31375.4]
  wire [7:0] _T_57542; // @[Mux.scala 19:72:@31382.4]
  wire [7:0] _T_57549; // @[Mux.scala 19:72:@31389.4]
  wire [15:0] _T_57550; // @[Mux.scala 19:72:@31390.4]
  wire [15:0] _T_57552; // @[Mux.scala 19:72:@31391.4]
  wire [7:0] _T_57559; // @[Mux.scala 19:72:@31398.4]
  wire [7:0] _T_57566; // @[Mux.scala 19:72:@31405.4]
  wire [15:0] _T_57567; // @[Mux.scala 19:72:@31406.4]
  wire [15:0] _T_57569; // @[Mux.scala 19:72:@31407.4]
  wire [7:0] _T_57576; // @[Mux.scala 19:72:@31414.4]
  wire [7:0] _T_57583; // @[Mux.scala 19:72:@31421.4]
  wire [15:0] _T_57584; // @[Mux.scala 19:72:@31422.4]
  wire [15:0] _T_57586; // @[Mux.scala 19:72:@31423.4]
  wire [7:0] _T_57593; // @[Mux.scala 19:72:@31430.4]
  wire [7:0] _T_57600; // @[Mux.scala 19:72:@31437.4]
  wire [15:0] _T_57601; // @[Mux.scala 19:72:@31438.4]
  wire [15:0] _T_57603; // @[Mux.scala 19:72:@31439.4]
  wire [15:0] _T_57618; // @[Mux.scala 19:72:@31454.4]
  wire [15:0] _T_57620; // @[Mux.scala 19:72:@31455.4]
  wire [15:0] _T_57635; // @[Mux.scala 19:72:@31470.4]
  wire [15:0] _T_57637; // @[Mux.scala 19:72:@31471.4]
  wire [15:0] _T_57652; // @[Mux.scala 19:72:@31486.4]
  wire [15:0] _T_57654; // @[Mux.scala 19:72:@31487.4]
  wire [15:0] _T_57669; // @[Mux.scala 19:72:@31502.4]
  wire [15:0] _T_57671; // @[Mux.scala 19:72:@31503.4]
  wire [15:0] _T_57686; // @[Mux.scala 19:72:@31518.4]
  wire [15:0] _T_57688; // @[Mux.scala 19:72:@31519.4]
  wire [15:0] _T_57703; // @[Mux.scala 19:72:@31534.4]
  wire [15:0] _T_57705; // @[Mux.scala 19:72:@31535.4]
  wire [15:0] _T_57720; // @[Mux.scala 19:72:@31550.4]
  wire [15:0] _T_57722; // @[Mux.scala 19:72:@31551.4]
  wire [15:0] _T_57737; // @[Mux.scala 19:72:@31566.4]
  wire [15:0] _T_57739; // @[Mux.scala 19:72:@31567.4]
  wire [15:0] _T_57740; // @[Mux.scala 19:72:@31568.4]
  wire [15:0] _T_57741; // @[Mux.scala 19:72:@31569.4]
  wire [15:0] _T_57742; // @[Mux.scala 19:72:@31570.4]
  wire [15:0] _T_57743; // @[Mux.scala 19:72:@31571.4]
  wire [15:0] _T_57744; // @[Mux.scala 19:72:@31572.4]
  wire [15:0] _T_57745; // @[Mux.scala 19:72:@31573.4]
  wire [15:0] _T_57746; // @[Mux.scala 19:72:@31574.4]
  wire [15:0] _T_57747; // @[Mux.scala 19:72:@31575.4]
  wire [15:0] _T_57748; // @[Mux.scala 19:72:@31576.4]
  wire [15:0] _T_57749; // @[Mux.scala 19:72:@31577.4]
  wire [15:0] _T_57750; // @[Mux.scala 19:72:@31578.4]
  wire [15:0] _T_57751; // @[Mux.scala 19:72:@31579.4]
  wire [15:0] _T_57752; // @[Mux.scala 19:72:@31580.4]
  wire [15:0] _T_57753; // @[Mux.scala 19:72:@31581.4]
  wire [15:0] _T_57754; // @[Mux.scala 19:72:@31582.4]
  wire [7:0] _T_58332; // @[Mux.scala 19:72:@31932.4]
  wire [7:0] _T_58339; // @[Mux.scala 19:72:@31939.4]
  wire [15:0] _T_58340; // @[Mux.scala 19:72:@31940.4]
  wire [15:0] _T_58342; // @[Mux.scala 19:72:@31941.4]
  wire [7:0] _T_58349; // @[Mux.scala 19:72:@31948.4]
  wire [7:0] _T_58356; // @[Mux.scala 19:72:@31955.4]
  wire [15:0] _T_58357; // @[Mux.scala 19:72:@31956.4]
  wire [15:0] _T_58359; // @[Mux.scala 19:72:@31957.4]
  wire [7:0] _T_58366; // @[Mux.scala 19:72:@31964.4]
  wire [7:0] _T_58373; // @[Mux.scala 19:72:@31971.4]
  wire [15:0] _T_58374; // @[Mux.scala 19:72:@31972.4]
  wire [15:0] _T_58376; // @[Mux.scala 19:72:@31973.4]
  wire [7:0] _T_58383; // @[Mux.scala 19:72:@31980.4]
  wire [7:0] _T_58390; // @[Mux.scala 19:72:@31987.4]
  wire [15:0] _T_58391; // @[Mux.scala 19:72:@31988.4]
  wire [15:0] _T_58393; // @[Mux.scala 19:72:@31989.4]
  wire [7:0] _T_58400; // @[Mux.scala 19:72:@31996.4]
  wire [7:0] _T_58407; // @[Mux.scala 19:72:@32003.4]
  wire [15:0] _T_58408; // @[Mux.scala 19:72:@32004.4]
  wire [15:0] _T_58410; // @[Mux.scala 19:72:@32005.4]
  wire [7:0] _T_58417; // @[Mux.scala 19:72:@32012.4]
  wire [7:0] _T_58424; // @[Mux.scala 19:72:@32019.4]
  wire [15:0] _T_58425; // @[Mux.scala 19:72:@32020.4]
  wire [15:0] _T_58427; // @[Mux.scala 19:72:@32021.4]
  wire [7:0] _T_58434; // @[Mux.scala 19:72:@32028.4]
  wire [7:0] _T_58441; // @[Mux.scala 19:72:@32035.4]
  wire [15:0] _T_58442; // @[Mux.scala 19:72:@32036.4]
  wire [15:0] _T_58444; // @[Mux.scala 19:72:@32037.4]
  wire [7:0] _T_58451; // @[Mux.scala 19:72:@32044.4]
  wire [7:0] _T_58458; // @[Mux.scala 19:72:@32051.4]
  wire [15:0] _T_58459; // @[Mux.scala 19:72:@32052.4]
  wire [15:0] _T_58461; // @[Mux.scala 19:72:@32053.4]
  wire [15:0] _T_58476; // @[Mux.scala 19:72:@32068.4]
  wire [15:0] _T_58478; // @[Mux.scala 19:72:@32069.4]
  wire [15:0] _T_58493; // @[Mux.scala 19:72:@32084.4]
  wire [15:0] _T_58495; // @[Mux.scala 19:72:@32085.4]
  wire [15:0] _T_58510; // @[Mux.scala 19:72:@32100.4]
  wire [15:0] _T_58512; // @[Mux.scala 19:72:@32101.4]
  wire [15:0] _T_58527; // @[Mux.scala 19:72:@32116.4]
  wire [15:0] _T_58529; // @[Mux.scala 19:72:@32117.4]
  wire [15:0] _T_58544; // @[Mux.scala 19:72:@32132.4]
  wire [15:0] _T_58546; // @[Mux.scala 19:72:@32133.4]
  wire [15:0] _T_58561; // @[Mux.scala 19:72:@32148.4]
  wire [15:0] _T_58563; // @[Mux.scala 19:72:@32149.4]
  wire [15:0] _T_58578; // @[Mux.scala 19:72:@32164.4]
  wire [15:0] _T_58580; // @[Mux.scala 19:72:@32165.4]
  wire [15:0] _T_58595; // @[Mux.scala 19:72:@32180.4]
  wire [15:0] _T_58597; // @[Mux.scala 19:72:@32181.4]
  wire [15:0] _T_58598; // @[Mux.scala 19:72:@32182.4]
  wire [15:0] _T_58599; // @[Mux.scala 19:72:@32183.4]
  wire [15:0] _T_58600; // @[Mux.scala 19:72:@32184.4]
  wire [15:0] _T_58601; // @[Mux.scala 19:72:@32185.4]
  wire [15:0] _T_58602; // @[Mux.scala 19:72:@32186.4]
  wire [15:0] _T_58603; // @[Mux.scala 19:72:@32187.4]
  wire [15:0] _T_58604; // @[Mux.scala 19:72:@32188.4]
  wire [15:0] _T_58605; // @[Mux.scala 19:72:@32189.4]
  wire [15:0] _T_58606; // @[Mux.scala 19:72:@32190.4]
  wire [15:0] _T_58607; // @[Mux.scala 19:72:@32191.4]
  wire [15:0] _T_58608; // @[Mux.scala 19:72:@32192.4]
  wire [15:0] _T_58609; // @[Mux.scala 19:72:@32193.4]
  wire [15:0] _T_58610; // @[Mux.scala 19:72:@32194.4]
  wire [15:0] _T_58611; // @[Mux.scala 19:72:@32195.4]
  wire [15:0] _T_58612; // @[Mux.scala 19:72:@32196.4]
  wire [7:0] _T_59190; // @[Mux.scala 19:72:@32546.4]
  wire [7:0] _T_59197; // @[Mux.scala 19:72:@32553.4]
  wire [15:0] _T_59198; // @[Mux.scala 19:72:@32554.4]
  wire [15:0] _T_59200; // @[Mux.scala 19:72:@32555.4]
  wire [7:0] _T_59207; // @[Mux.scala 19:72:@32562.4]
  wire [7:0] _T_59214; // @[Mux.scala 19:72:@32569.4]
  wire [15:0] _T_59215; // @[Mux.scala 19:72:@32570.4]
  wire [15:0] _T_59217; // @[Mux.scala 19:72:@32571.4]
  wire [7:0] _T_59224; // @[Mux.scala 19:72:@32578.4]
  wire [7:0] _T_59231; // @[Mux.scala 19:72:@32585.4]
  wire [15:0] _T_59232; // @[Mux.scala 19:72:@32586.4]
  wire [15:0] _T_59234; // @[Mux.scala 19:72:@32587.4]
  wire [7:0] _T_59241; // @[Mux.scala 19:72:@32594.4]
  wire [7:0] _T_59248; // @[Mux.scala 19:72:@32601.4]
  wire [15:0] _T_59249; // @[Mux.scala 19:72:@32602.4]
  wire [15:0] _T_59251; // @[Mux.scala 19:72:@32603.4]
  wire [7:0] _T_59258; // @[Mux.scala 19:72:@32610.4]
  wire [7:0] _T_59265; // @[Mux.scala 19:72:@32617.4]
  wire [15:0] _T_59266; // @[Mux.scala 19:72:@32618.4]
  wire [15:0] _T_59268; // @[Mux.scala 19:72:@32619.4]
  wire [7:0] _T_59275; // @[Mux.scala 19:72:@32626.4]
  wire [7:0] _T_59282; // @[Mux.scala 19:72:@32633.4]
  wire [15:0] _T_59283; // @[Mux.scala 19:72:@32634.4]
  wire [15:0] _T_59285; // @[Mux.scala 19:72:@32635.4]
  wire [7:0] _T_59292; // @[Mux.scala 19:72:@32642.4]
  wire [7:0] _T_59299; // @[Mux.scala 19:72:@32649.4]
  wire [15:0] _T_59300; // @[Mux.scala 19:72:@32650.4]
  wire [15:0] _T_59302; // @[Mux.scala 19:72:@32651.4]
  wire [7:0] _T_59309; // @[Mux.scala 19:72:@32658.4]
  wire [7:0] _T_59316; // @[Mux.scala 19:72:@32665.4]
  wire [15:0] _T_59317; // @[Mux.scala 19:72:@32666.4]
  wire [15:0] _T_59319; // @[Mux.scala 19:72:@32667.4]
  wire [15:0] _T_59334; // @[Mux.scala 19:72:@32682.4]
  wire [15:0] _T_59336; // @[Mux.scala 19:72:@32683.4]
  wire [15:0] _T_59351; // @[Mux.scala 19:72:@32698.4]
  wire [15:0] _T_59353; // @[Mux.scala 19:72:@32699.4]
  wire [15:0] _T_59368; // @[Mux.scala 19:72:@32714.4]
  wire [15:0] _T_59370; // @[Mux.scala 19:72:@32715.4]
  wire [15:0] _T_59385; // @[Mux.scala 19:72:@32730.4]
  wire [15:0] _T_59387; // @[Mux.scala 19:72:@32731.4]
  wire [15:0] _T_59402; // @[Mux.scala 19:72:@32746.4]
  wire [15:0] _T_59404; // @[Mux.scala 19:72:@32747.4]
  wire [15:0] _T_59419; // @[Mux.scala 19:72:@32762.4]
  wire [15:0] _T_59421; // @[Mux.scala 19:72:@32763.4]
  wire [15:0] _T_59436; // @[Mux.scala 19:72:@32778.4]
  wire [15:0] _T_59438; // @[Mux.scala 19:72:@32779.4]
  wire [15:0] _T_59453; // @[Mux.scala 19:72:@32794.4]
  wire [15:0] _T_59455; // @[Mux.scala 19:72:@32795.4]
  wire [15:0] _T_59456; // @[Mux.scala 19:72:@32796.4]
  wire [15:0] _T_59457; // @[Mux.scala 19:72:@32797.4]
  wire [15:0] _T_59458; // @[Mux.scala 19:72:@32798.4]
  wire [15:0] _T_59459; // @[Mux.scala 19:72:@32799.4]
  wire [15:0] _T_59460; // @[Mux.scala 19:72:@32800.4]
  wire [15:0] _T_59461; // @[Mux.scala 19:72:@32801.4]
  wire [15:0] _T_59462; // @[Mux.scala 19:72:@32802.4]
  wire [15:0] _T_59463; // @[Mux.scala 19:72:@32803.4]
  wire [15:0] _T_59464; // @[Mux.scala 19:72:@32804.4]
  wire [15:0] _T_59465; // @[Mux.scala 19:72:@32805.4]
  wire [15:0] _T_59466; // @[Mux.scala 19:72:@32806.4]
  wire [15:0] _T_59467; // @[Mux.scala 19:72:@32807.4]
  wire [15:0] _T_59468; // @[Mux.scala 19:72:@32808.4]
  wire [15:0] _T_59469; // @[Mux.scala 19:72:@32809.4]
  wire [15:0] _T_59470; // @[Mux.scala 19:72:@32810.4]
  wire [7:0] _T_60048; // @[Mux.scala 19:72:@33160.4]
  wire [7:0] _T_60055; // @[Mux.scala 19:72:@33167.4]
  wire [15:0] _T_60056; // @[Mux.scala 19:72:@33168.4]
  wire [15:0] _T_60058; // @[Mux.scala 19:72:@33169.4]
  wire [7:0] _T_60065; // @[Mux.scala 19:72:@33176.4]
  wire [7:0] _T_60072; // @[Mux.scala 19:72:@33183.4]
  wire [15:0] _T_60073; // @[Mux.scala 19:72:@33184.4]
  wire [15:0] _T_60075; // @[Mux.scala 19:72:@33185.4]
  wire [7:0] _T_60082; // @[Mux.scala 19:72:@33192.4]
  wire [7:0] _T_60089; // @[Mux.scala 19:72:@33199.4]
  wire [15:0] _T_60090; // @[Mux.scala 19:72:@33200.4]
  wire [15:0] _T_60092; // @[Mux.scala 19:72:@33201.4]
  wire [7:0] _T_60099; // @[Mux.scala 19:72:@33208.4]
  wire [7:0] _T_60106; // @[Mux.scala 19:72:@33215.4]
  wire [15:0] _T_60107; // @[Mux.scala 19:72:@33216.4]
  wire [15:0] _T_60109; // @[Mux.scala 19:72:@33217.4]
  wire [7:0] _T_60116; // @[Mux.scala 19:72:@33224.4]
  wire [7:0] _T_60123; // @[Mux.scala 19:72:@33231.4]
  wire [15:0] _T_60124; // @[Mux.scala 19:72:@33232.4]
  wire [15:0] _T_60126; // @[Mux.scala 19:72:@33233.4]
  wire [7:0] _T_60133; // @[Mux.scala 19:72:@33240.4]
  wire [7:0] _T_60140; // @[Mux.scala 19:72:@33247.4]
  wire [15:0] _T_60141; // @[Mux.scala 19:72:@33248.4]
  wire [15:0] _T_60143; // @[Mux.scala 19:72:@33249.4]
  wire [7:0] _T_60150; // @[Mux.scala 19:72:@33256.4]
  wire [7:0] _T_60157; // @[Mux.scala 19:72:@33263.4]
  wire [15:0] _T_60158; // @[Mux.scala 19:72:@33264.4]
  wire [15:0] _T_60160; // @[Mux.scala 19:72:@33265.4]
  wire [7:0] _T_60167; // @[Mux.scala 19:72:@33272.4]
  wire [7:0] _T_60174; // @[Mux.scala 19:72:@33279.4]
  wire [15:0] _T_60175; // @[Mux.scala 19:72:@33280.4]
  wire [15:0] _T_60177; // @[Mux.scala 19:72:@33281.4]
  wire [15:0] _T_60192; // @[Mux.scala 19:72:@33296.4]
  wire [15:0] _T_60194; // @[Mux.scala 19:72:@33297.4]
  wire [15:0] _T_60209; // @[Mux.scala 19:72:@33312.4]
  wire [15:0] _T_60211; // @[Mux.scala 19:72:@33313.4]
  wire [15:0] _T_60226; // @[Mux.scala 19:72:@33328.4]
  wire [15:0] _T_60228; // @[Mux.scala 19:72:@33329.4]
  wire [15:0] _T_60243; // @[Mux.scala 19:72:@33344.4]
  wire [15:0] _T_60245; // @[Mux.scala 19:72:@33345.4]
  wire [15:0] _T_60260; // @[Mux.scala 19:72:@33360.4]
  wire [15:0] _T_60262; // @[Mux.scala 19:72:@33361.4]
  wire [15:0] _T_60277; // @[Mux.scala 19:72:@33376.4]
  wire [15:0] _T_60279; // @[Mux.scala 19:72:@33377.4]
  wire [15:0] _T_60294; // @[Mux.scala 19:72:@33392.4]
  wire [15:0] _T_60296; // @[Mux.scala 19:72:@33393.4]
  wire [15:0] _T_60311; // @[Mux.scala 19:72:@33408.4]
  wire [15:0] _T_60313; // @[Mux.scala 19:72:@33409.4]
  wire [15:0] _T_60314; // @[Mux.scala 19:72:@33410.4]
  wire [15:0] _T_60315; // @[Mux.scala 19:72:@33411.4]
  wire [15:0] _T_60316; // @[Mux.scala 19:72:@33412.4]
  wire [15:0] _T_60317; // @[Mux.scala 19:72:@33413.4]
  wire [15:0] _T_60318; // @[Mux.scala 19:72:@33414.4]
  wire [15:0] _T_60319; // @[Mux.scala 19:72:@33415.4]
  wire [15:0] _T_60320; // @[Mux.scala 19:72:@33416.4]
  wire [15:0] _T_60321; // @[Mux.scala 19:72:@33417.4]
  wire [15:0] _T_60322; // @[Mux.scala 19:72:@33418.4]
  wire [15:0] _T_60323; // @[Mux.scala 19:72:@33419.4]
  wire [15:0] _T_60324; // @[Mux.scala 19:72:@33420.4]
  wire [15:0] _T_60325; // @[Mux.scala 19:72:@33421.4]
  wire [15:0] _T_60326; // @[Mux.scala 19:72:@33422.4]
  wire [15:0] _T_60327; // @[Mux.scala 19:72:@33423.4]
  wire [15:0] _T_60328; // @[Mux.scala 19:72:@33424.4]
  wire [7:0] _T_60906; // @[Mux.scala 19:72:@33774.4]
  wire [7:0] _T_60913; // @[Mux.scala 19:72:@33781.4]
  wire [15:0] _T_60914; // @[Mux.scala 19:72:@33782.4]
  wire [15:0] _T_60916; // @[Mux.scala 19:72:@33783.4]
  wire [7:0] _T_60923; // @[Mux.scala 19:72:@33790.4]
  wire [7:0] _T_60930; // @[Mux.scala 19:72:@33797.4]
  wire [15:0] _T_60931; // @[Mux.scala 19:72:@33798.4]
  wire [15:0] _T_60933; // @[Mux.scala 19:72:@33799.4]
  wire [7:0] _T_60940; // @[Mux.scala 19:72:@33806.4]
  wire [7:0] _T_60947; // @[Mux.scala 19:72:@33813.4]
  wire [15:0] _T_60948; // @[Mux.scala 19:72:@33814.4]
  wire [15:0] _T_60950; // @[Mux.scala 19:72:@33815.4]
  wire [7:0] _T_60957; // @[Mux.scala 19:72:@33822.4]
  wire [7:0] _T_60964; // @[Mux.scala 19:72:@33829.4]
  wire [15:0] _T_60965; // @[Mux.scala 19:72:@33830.4]
  wire [15:0] _T_60967; // @[Mux.scala 19:72:@33831.4]
  wire [7:0] _T_60974; // @[Mux.scala 19:72:@33838.4]
  wire [7:0] _T_60981; // @[Mux.scala 19:72:@33845.4]
  wire [15:0] _T_60982; // @[Mux.scala 19:72:@33846.4]
  wire [15:0] _T_60984; // @[Mux.scala 19:72:@33847.4]
  wire [7:0] _T_60991; // @[Mux.scala 19:72:@33854.4]
  wire [7:0] _T_60998; // @[Mux.scala 19:72:@33861.4]
  wire [15:0] _T_60999; // @[Mux.scala 19:72:@33862.4]
  wire [15:0] _T_61001; // @[Mux.scala 19:72:@33863.4]
  wire [7:0] _T_61008; // @[Mux.scala 19:72:@33870.4]
  wire [7:0] _T_61015; // @[Mux.scala 19:72:@33877.4]
  wire [15:0] _T_61016; // @[Mux.scala 19:72:@33878.4]
  wire [15:0] _T_61018; // @[Mux.scala 19:72:@33879.4]
  wire [7:0] _T_61025; // @[Mux.scala 19:72:@33886.4]
  wire [7:0] _T_61032; // @[Mux.scala 19:72:@33893.4]
  wire [15:0] _T_61033; // @[Mux.scala 19:72:@33894.4]
  wire [15:0] _T_61035; // @[Mux.scala 19:72:@33895.4]
  wire [15:0] _T_61050; // @[Mux.scala 19:72:@33910.4]
  wire [15:0] _T_61052; // @[Mux.scala 19:72:@33911.4]
  wire [15:0] _T_61067; // @[Mux.scala 19:72:@33926.4]
  wire [15:0] _T_61069; // @[Mux.scala 19:72:@33927.4]
  wire [15:0] _T_61084; // @[Mux.scala 19:72:@33942.4]
  wire [15:0] _T_61086; // @[Mux.scala 19:72:@33943.4]
  wire [15:0] _T_61101; // @[Mux.scala 19:72:@33958.4]
  wire [15:0] _T_61103; // @[Mux.scala 19:72:@33959.4]
  wire [15:0] _T_61118; // @[Mux.scala 19:72:@33974.4]
  wire [15:0] _T_61120; // @[Mux.scala 19:72:@33975.4]
  wire [15:0] _T_61135; // @[Mux.scala 19:72:@33990.4]
  wire [15:0] _T_61137; // @[Mux.scala 19:72:@33991.4]
  wire [15:0] _T_61152; // @[Mux.scala 19:72:@34006.4]
  wire [15:0] _T_61154; // @[Mux.scala 19:72:@34007.4]
  wire [15:0] _T_61169; // @[Mux.scala 19:72:@34022.4]
  wire [15:0] _T_61171; // @[Mux.scala 19:72:@34023.4]
  wire [15:0] _T_61172; // @[Mux.scala 19:72:@34024.4]
  wire [15:0] _T_61173; // @[Mux.scala 19:72:@34025.4]
  wire [15:0] _T_61174; // @[Mux.scala 19:72:@34026.4]
  wire [15:0] _T_61175; // @[Mux.scala 19:72:@34027.4]
  wire [15:0] _T_61176; // @[Mux.scala 19:72:@34028.4]
  wire [15:0] _T_61177; // @[Mux.scala 19:72:@34029.4]
  wire [15:0] _T_61178; // @[Mux.scala 19:72:@34030.4]
  wire [15:0] _T_61179; // @[Mux.scala 19:72:@34031.4]
  wire [15:0] _T_61180; // @[Mux.scala 19:72:@34032.4]
  wire [15:0] _T_61181; // @[Mux.scala 19:72:@34033.4]
  wire [15:0] _T_61182; // @[Mux.scala 19:72:@34034.4]
  wire [15:0] _T_61183; // @[Mux.scala 19:72:@34035.4]
  wire [15:0] _T_61184; // @[Mux.scala 19:72:@34036.4]
  wire [15:0] _T_61185; // @[Mux.scala 19:72:@34037.4]
  wire [15:0] _T_61186; // @[Mux.scala 19:72:@34038.4]
  wire [7:0] _T_61764; // @[Mux.scala 19:72:@34388.4]
  wire [7:0] _T_61771; // @[Mux.scala 19:72:@34395.4]
  wire [15:0] _T_61772; // @[Mux.scala 19:72:@34396.4]
  wire [15:0] _T_61774; // @[Mux.scala 19:72:@34397.4]
  wire [7:0] _T_61781; // @[Mux.scala 19:72:@34404.4]
  wire [7:0] _T_61788; // @[Mux.scala 19:72:@34411.4]
  wire [15:0] _T_61789; // @[Mux.scala 19:72:@34412.4]
  wire [15:0] _T_61791; // @[Mux.scala 19:72:@34413.4]
  wire [7:0] _T_61798; // @[Mux.scala 19:72:@34420.4]
  wire [7:0] _T_61805; // @[Mux.scala 19:72:@34427.4]
  wire [15:0] _T_61806; // @[Mux.scala 19:72:@34428.4]
  wire [15:0] _T_61808; // @[Mux.scala 19:72:@34429.4]
  wire [7:0] _T_61815; // @[Mux.scala 19:72:@34436.4]
  wire [7:0] _T_61822; // @[Mux.scala 19:72:@34443.4]
  wire [15:0] _T_61823; // @[Mux.scala 19:72:@34444.4]
  wire [15:0] _T_61825; // @[Mux.scala 19:72:@34445.4]
  wire [7:0] _T_61832; // @[Mux.scala 19:72:@34452.4]
  wire [7:0] _T_61839; // @[Mux.scala 19:72:@34459.4]
  wire [15:0] _T_61840; // @[Mux.scala 19:72:@34460.4]
  wire [15:0] _T_61842; // @[Mux.scala 19:72:@34461.4]
  wire [7:0] _T_61849; // @[Mux.scala 19:72:@34468.4]
  wire [7:0] _T_61856; // @[Mux.scala 19:72:@34475.4]
  wire [15:0] _T_61857; // @[Mux.scala 19:72:@34476.4]
  wire [15:0] _T_61859; // @[Mux.scala 19:72:@34477.4]
  wire [7:0] _T_61866; // @[Mux.scala 19:72:@34484.4]
  wire [7:0] _T_61873; // @[Mux.scala 19:72:@34491.4]
  wire [15:0] _T_61874; // @[Mux.scala 19:72:@34492.4]
  wire [15:0] _T_61876; // @[Mux.scala 19:72:@34493.4]
  wire [7:0] _T_61883; // @[Mux.scala 19:72:@34500.4]
  wire [7:0] _T_61890; // @[Mux.scala 19:72:@34507.4]
  wire [15:0] _T_61891; // @[Mux.scala 19:72:@34508.4]
  wire [15:0] _T_61893; // @[Mux.scala 19:72:@34509.4]
  wire [15:0] _T_61908; // @[Mux.scala 19:72:@34524.4]
  wire [15:0] _T_61910; // @[Mux.scala 19:72:@34525.4]
  wire [15:0] _T_61925; // @[Mux.scala 19:72:@34540.4]
  wire [15:0] _T_61927; // @[Mux.scala 19:72:@34541.4]
  wire [15:0] _T_61942; // @[Mux.scala 19:72:@34556.4]
  wire [15:0] _T_61944; // @[Mux.scala 19:72:@34557.4]
  wire [15:0] _T_61959; // @[Mux.scala 19:72:@34572.4]
  wire [15:0] _T_61961; // @[Mux.scala 19:72:@34573.4]
  wire [15:0] _T_61976; // @[Mux.scala 19:72:@34588.4]
  wire [15:0] _T_61978; // @[Mux.scala 19:72:@34589.4]
  wire [15:0] _T_61993; // @[Mux.scala 19:72:@34604.4]
  wire [15:0] _T_61995; // @[Mux.scala 19:72:@34605.4]
  wire [15:0] _T_62010; // @[Mux.scala 19:72:@34620.4]
  wire [15:0] _T_62012; // @[Mux.scala 19:72:@34621.4]
  wire [15:0] _T_62027; // @[Mux.scala 19:72:@34636.4]
  wire [15:0] _T_62029; // @[Mux.scala 19:72:@34637.4]
  wire [15:0] _T_62030; // @[Mux.scala 19:72:@34638.4]
  wire [15:0] _T_62031; // @[Mux.scala 19:72:@34639.4]
  wire [15:0] _T_62032; // @[Mux.scala 19:72:@34640.4]
  wire [15:0] _T_62033; // @[Mux.scala 19:72:@34641.4]
  wire [15:0] _T_62034; // @[Mux.scala 19:72:@34642.4]
  wire [15:0] _T_62035; // @[Mux.scala 19:72:@34643.4]
  wire [15:0] _T_62036; // @[Mux.scala 19:72:@34644.4]
  wire [15:0] _T_62037; // @[Mux.scala 19:72:@34645.4]
  wire [15:0] _T_62038; // @[Mux.scala 19:72:@34646.4]
  wire [15:0] _T_62039; // @[Mux.scala 19:72:@34647.4]
  wire [15:0] _T_62040; // @[Mux.scala 19:72:@34648.4]
  wire [15:0] _T_62041; // @[Mux.scala 19:72:@34649.4]
  wire [15:0] _T_62042; // @[Mux.scala 19:72:@34650.4]
  wire [15:0] _T_62043; // @[Mux.scala 19:72:@34651.4]
  wire [15:0] _T_62044; // @[Mux.scala 19:72:@34652.4]
  wire [7:0] _T_62622; // @[Mux.scala 19:72:@35002.4]
  wire [7:0] _T_62629; // @[Mux.scala 19:72:@35009.4]
  wire [15:0] _T_62630; // @[Mux.scala 19:72:@35010.4]
  wire [15:0] _T_62632; // @[Mux.scala 19:72:@35011.4]
  wire [7:0] _T_62639; // @[Mux.scala 19:72:@35018.4]
  wire [7:0] _T_62646; // @[Mux.scala 19:72:@35025.4]
  wire [15:0] _T_62647; // @[Mux.scala 19:72:@35026.4]
  wire [15:0] _T_62649; // @[Mux.scala 19:72:@35027.4]
  wire [7:0] _T_62656; // @[Mux.scala 19:72:@35034.4]
  wire [7:0] _T_62663; // @[Mux.scala 19:72:@35041.4]
  wire [15:0] _T_62664; // @[Mux.scala 19:72:@35042.4]
  wire [15:0] _T_62666; // @[Mux.scala 19:72:@35043.4]
  wire [7:0] _T_62673; // @[Mux.scala 19:72:@35050.4]
  wire [7:0] _T_62680; // @[Mux.scala 19:72:@35057.4]
  wire [15:0] _T_62681; // @[Mux.scala 19:72:@35058.4]
  wire [15:0] _T_62683; // @[Mux.scala 19:72:@35059.4]
  wire [7:0] _T_62690; // @[Mux.scala 19:72:@35066.4]
  wire [7:0] _T_62697; // @[Mux.scala 19:72:@35073.4]
  wire [15:0] _T_62698; // @[Mux.scala 19:72:@35074.4]
  wire [15:0] _T_62700; // @[Mux.scala 19:72:@35075.4]
  wire [7:0] _T_62707; // @[Mux.scala 19:72:@35082.4]
  wire [7:0] _T_62714; // @[Mux.scala 19:72:@35089.4]
  wire [15:0] _T_62715; // @[Mux.scala 19:72:@35090.4]
  wire [15:0] _T_62717; // @[Mux.scala 19:72:@35091.4]
  wire [7:0] _T_62724; // @[Mux.scala 19:72:@35098.4]
  wire [7:0] _T_62731; // @[Mux.scala 19:72:@35105.4]
  wire [15:0] _T_62732; // @[Mux.scala 19:72:@35106.4]
  wire [15:0] _T_62734; // @[Mux.scala 19:72:@35107.4]
  wire [7:0] _T_62741; // @[Mux.scala 19:72:@35114.4]
  wire [7:0] _T_62748; // @[Mux.scala 19:72:@35121.4]
  wire [15:0] _T_62749; // @[Mux.scala 19:72:@35122.4]
  wire [15:0] _T_62751; // @[Mux.scala 19:72:@35123.4]
  wire [15:0] _T_62766; // @[Mux.scala 19:72:@35138.4]
  wire [15:0] _T_62768; // @[Mux.scala 19:72:@35139.4]
  wire [15:0] _T_62783; // @[Mux.scala 19:72:@35154.4]
  wire [15:0] _T_62785; // @[Mux.scala 19:72:@35155.4]
  wire [15:0] _T_62800; // @[Mux.scala 19:72:@35170.4]
  wire [15:0] _T_62802; // @[Mux.scala 19:72:@35171.4]
  wire [15:0] _T_62817; // @[Mux.scala 19:72:@35186.4]
  wire [15:0] _T_62819; // @[Mux.scala 19:72:@35187.4]
  wire [15:0] _T_62834; // @[Mux.scala 19:72:@35202.4]
  wire [15:0] _T_62836; // @[Mux.scala 19:72:@35203.4]
  wire [15:0] _T_62851; // @[Mux.scala 19:72:@35218.4]
  wire [15:0] _T_62853; // @[Mux.scala 19:72:@35219.4]
  wire [15:0] _T_62868; // @[Mux.scala 19:72:@35234.4]
  wire [15:0] _T_62870; // @[Mux.scala 19:72:@35235.4]
  wire [15:0] _T_62885; // @[Mux.scala 19:72:@35250.4]
  wire [15:0] _T_62887; // @[Mux.scala 19:72:@35251.4]
  wire [15:0] _T_62888; // @[Mux.scala 19:72:@35252.4]
  wire [15:0] _T_62889; // @[Mux.scala 19:72:@35253.4]
  wire [15:0] _T_62890; // @[Mux.scala 19:72:@35254.4]
  wire [15:0] _T_62891; // @[Mux.scala 19:72:@35255.4]
  wire [15:0] _T_62892; // @[Mux.scala 19:72:@35256.4]
  wire [15:0] _T_62893; // @[Mux.scala 19:72:@35257.4]
  wire [15:0] _T_62894; // @[Mux.scala 19:72:@35258.4]
  wire [15:0] _T_62895; // @[Mux.scala 19:72:@35259.4]
  wire [15:0] _T_62896; // @[Mux.scala 19:72:@35260.4]
  wire [15:0] _T_62897; // @[Mux.scala 19:72:@35261.4]
  wire [15:0] _T_62898; // @[Mux.scala 19:72:@35262.4]
  wire [15:0] _T_62899; // @[Mux.scala 19:72:@35263.4]
  wire [15:0] _T_62900; // @[Mux.scala 19:72:@35264.4]
  wire [15:0] _T_62901; // @[Mux.scala 19:72:@35265.4]
  wire [15:0] _T_62902; // @[Mux.scala 19:72:@35266.4]
  wire [7:0] _T_63480; // @[Mux.scala 19:72:@35616.4]
  wire [7:0] _T_63487; // @[Mux.scala 19:72:@35623.4]
  wire [15:0] _T_63488; // @[Mux.scala 19:72:@35624.4]
  wire [15:0] _T_63490; // @[Mux.scala 19:72:@35625.4]
  wire [7:0] _T_63497; // @[Mux.scala 19:72:@35632.4]
  wire [7:0] _T_63504; // @[Mux.scala 19:72:@35639.4]
  wire [15:0] _T_63505; // @[Mux.scala 19:72:@35640.4]
  wire [15:0] _T_63507; // @[Mux.scala 19:72:@35641.4]
  wire [7:0] _T_63514; // @[Mux.scala 19:72:@35648.4]
  wire [7:0] _T_63521; // @[Mux.scala 19:72:@35655.4]
  wire [15:0] _T_63522; // @[Mux.scala 19:72:@35656.4]
  wire [15:0] _T_63524; // @[Mux.scala 19:72:@35657.4]
  wire [7:0] _T_63531; // @[Mux.scala 19:72:@35664.4]
  wire [7:0] _T_63538; // @[Mux.scala 19:72:@35671.4]
  wire [15:0] _T_63539; // @[Mux.scala 19:72:@35672.4]
  wire [15:0] _T_63541; // @[Mux.scala 19:72:@35673.4]
  wire [7:0] _T_63548; // @[Mux.scala 19:72:@35680.4]
  wire [7:0] _T_63555; // @[Mux.scala 19:72:@35687.4]
  wire [15:0] _T_63556; // @[Mux.scala 19:72:@35688.4]
  wire [15:0] _T_63558; // @[Mux.scala 19:72:@35689.4]
  wire [7:0] _T_63565; // @[Mux.scala 19:72:@35696.4]
  wire [7:0] _T_63572; // @[Mux.scala 19:72:@35703.4]
  wire [15:0] _T_63573; // @[Mux.scala 19:72:@35704.4]
  wire [15:0] _T_63575; // @[Mux.scala 19:72:@35705.4]
  wire [7:0] _T_63582; // @[Mux.scala 19:72:@35712.4]
  wire [7:0] _T_63589; // @[Mux.scala 19:72:@35719.4]
  wire [15:0] _T_63590; // @[Mux.scala 19:72:@35720.4]
  wire [15:0] _T_63592; // @[Mux.scala 19:72:@35721.4]
  wire [7:0] _T_63599; // @[Mux.scala 19:72:@35728.4]
  wire [7:0] _T_63606; // @[Mux.scala 19:72:@35735.4]
  wire [15:0] _T_63607; // @[Mux.scala 19:72:@35736.4]
  wire [15:0] _T_63609; // @[Mux.scala 19:72:@35737.4]
  wire [15:0] _T_63624; // @[Mux.scala 19:72:@35752.4]
  wire [15:0] _T_63626; // @[Mux.scala 19:72:@35753.4]
  wire [15:0] _T_63641; // @[Mux.scala 19:72:@35768.4]
  wire [15:0] _T_63643; // @[Mux.scala 19:72:@35769.4]
  wire [15:0] _T_63658; // @[Mux.scala 19:72:@35784.4]
  wire [15:0] _T_63660; // @[Mux.scala 19:72:@35785.4]
  wire [15:0] _T_63675; // @[Mux.scala 19:72:@35800.4]
  wire [15:0] _T_63677; // @[Mux.scala 19:72:@35801.4]
  wire [15:0] _T_63692; // @[Mux.scala 19:72:@35816.4]
  wire [15:0] _T_63694; // @[Mux.scala 19:72:@35817.4]
  wire [15:0] _T_63709; // @[Mux.scala 19:72:@35832.4]
  wire [15:0] _T_63711; // @[Mux.scala 19:72:@35833.4]
  wire [15:0] _T_63726; // @[Mux.scala 19:72:@35848.4]
  wire [15:0] _T_63728; // @[Mux.scala 19:72:@35849.4]
  wire [15:0] _T_63743; // @[Mux.scala 19:72:@35864.4]
  wire [15:0] _T_63745; // @[Mux.scala 19:72:@35865.4]
  wire [15:0] _T_63746; // @[Mux.scala 19:72:@35866.4]
  wire [15:0] _T_63747; // @[Mux.scala 19:72:@35867.4]
  wire [15:0] _T_63748; // @[Mux.scala 19:72:@35868.4]
  wire [15:0] _T_63749; // @[Mux.scala 19:72:@35869.4]
  wire [15:0] _T_63750; // @[Mux.scala 19:72:@35870.4]
  wire [15:0] _T_63751; // @[Mux.scala 19:72:@35871.4]
  wire [15:0] _T_63752; // @[Mux.scala 19:72:@35872.4]
  wire [15:0] _T_63753; // @[Mux.scala 19:72:@35873.4]
  wire [15:0] _T_63754; // @[Mux.scala 19:72:@35874.4]
  wire [15:0] _T_63755; // @[Mux.scala 19:72:@35875.4]
  wire [15:0] _T_63756; // @[Mux.scala 19:72:@35876.4]
  wire [15:0] _T_63757; // @[Mux.scala 19:72:@35877.4]
  wire [15:0] _T_63758; // @[Mux.scala 19:72:@35878.4]
  wire [15:0] _T_63759; // @[Mux.scala 19:72:@35879.4]
  wire [15:0] _T_63760; // @[Mux.scala 19:72:@35880.4]
  wire [7:0] _T_64338; // @[Mux.scala 19:72:@36230.4]
  wire [7:0] _T_64345; // @[Mux.scala 19:72:@36237.4]
  wire [15:0] _T_64346; // @[Mux.scala 19:72:@36238.4]
  wire [15:0] _T_64348; // @[Mux.scala 19:72:@36239.4]
  wire [7:0] _T_64355; // @[Mux.scala 19:72:@36246.4]
  wire [7:0] _T_64362; // @[Mux.scala 19:72:@36253.4]
  wire [15:0] _T_64363; // @[Mux.scala 19:72:@36254.4]
  wire [15:0] _T_64365; // @[Mux.scala 19:72:@36255.4]
  wire [7:0] _T_64372; // @[Mux.scala 19:72:@36262.4]
  wire [7:0] _T_64379; // @[Mux.scala 19:72:@36269.4]
  wire [15:0] _T_64380; // @[Mux.scala 19:72:@36270.4]
  wire [15:0] _T_64382; // @[Mux.scala 19:72:@36271.4]
  wire [7:0] _T_64389; // @[Mux.scala 19:72:@36278.4]
  wire [7:0] _T_64396; // @[Mux.scala 19:72:@36285.4]
  wire [15:0] _T_64397; // @[Mux.scala 19:72:@36286.4]
  wire [15:0] _T_64399; // @[Mux.scala 19:72:@36287.4]
  wire [7:0] _T_64406; // @[Mux.scala 19:72:@36294.4]
  wire [7:0] _T_64413; // @[Mux.scala 19:72:@36301.4]
  wire [15:0] _T_64414; // @[Mux.scala 19:72:@36302.4]
  wire [15:0] _T_64416; // @[Mux.scala 19:72:@36303.4]
  wire [7:0] _T_64423; // @[Mux.scala 19:72:@36310.4]
  wire [7:0] _T_64430; // @[Mux.scala 19:72:@36317.4]
  wire [15:0] _T_64431; // @[Mux.scala 19:72:@36318.4]
  wire [15:0] _T_64433; // @[Mux.scala 19:72:@36319.4]
  wire [7:0] _T_64440; // @[Mux.scala 19:72:@36326.4]
  wire [7:0] _T_64447; // @[Mux.scala 19:72:@36333.4]
  wire [15:0] _T_64448; // @[Mux.scala 19:72:@36334.4]
  wire [15:0] _T_64450; // @[Mux.scala 19:72:@36335.4]
  wire [7:0] _T_64457; // @[Mux.scala 19:72:@36342.4]
  wire [7:0] _T_64464; // @[Mux.scala 19:72:@36349.4]
  wire [15:0] _T_64465; // @[Mux.scala 19:72:@36350.4]
  wire [15:0] _T_64467; // @[Mux.scala 19:72:@36351.4]
  wire [15:0] _T_64482; // @[Mux.scala 19:72:@36366.4]
  wire [15:0] _T_64484; // @[Mux.scala 19:72:@36367.4]
  wire [15:0] _T_64499; // @[Mux.scala 19:72:@36382.4]
  wire [15:0] _T_64501; // @[Mux.scala 19:72:@36383.4]
  wire [15:0] _T_64516; // @[Mux.scala 19:72:@36398.4]
  wire [15:0] _T_64518; // @[Mux.scala 19:72:@36399.4]
  wire [15:0] _T_64533; // @[Mux.scala 19:72:@36414.4]
  wire [15:0] _T_64535; // @[Mux.scala 19:72:@36415.4]
  wire [15:0] _T_64550; // @[Mux.scala 19:72:@36430.4]
  wire [15:0] _T_64552; // @[Mux.scala 19:72:@36431.4]
  wire [15:0] _T_64567; // @[Mux.scala 19:72:@36446.4]
  wire [15:0] _T_64569; // @[Mux.scala 19:72:@36447.4]
  wire [15:0] _T_64584; // @[Mux.scala 19:72:@36462.4]
  wire [15:0] _T_64586; // @[Mux.scala 19:72:@36463.4]
  wire [15:0] _T_64601; // @[Mux.scala 19:72:@36478.4]
  wire [15:0] _T_64603; // @[Mux.scala 19:72:@36479.4]
  wire [15:0] _T_64604; // @[Mux.scala 19:72:@36480.4]
  wire [15:0] _T_64605; // @[Mux.scala 19:72:@36481.4]
  wire [15:0] _T_64606; // @[Mux.scala 19:72:@36482.4]
  wire [15:0] _T_64607; // @[Mux.scala 19:72:@36483.4]
  wire [15:0] _T_64608; // @[Mux.scala 19:72:@36484.4]
  wire [15:0] _T_64609; // @[Mux.scala 19:72:@36485.4]
  wire [15:0] _T_64610; // @[Mux.scala 19:72:@36486.4]
  wire [15:0] _T_64611; // @[Mux.scala 19:72:@36487.4]
  wire [15:0] _T_64612; // @[Mux.scala 19:72:@36488.4]
  wire [15:0] _T_64613; // @[Mux.scala 19:72:@36489.4]
  wire [15:0] _T_64614; // @[Mux.scala 19:72:@36490.4]
  wire [15:0] _T_64615; // @[Mux.scala 19:72:@36491.4]
  wire [15:0] _T_64616; // @[Mux.scala 19:72:@36492.4]
  wire [15:0] _T_64617; // @[Mux.scala 19:72:@36493.4]
  wire [15:0] _T_64618; // @[Mux.scala 19:72:@36494.4]
  wire [7:0] _T_65196; // @[Mux.scala 19:72:@36844.4]
  wire [7:0] _T_65203; // @[Mux.scala 19:72:@36851.4]
  wire [15:0] _T_65204; // @[Mux.scala 19:72:@36852.4]
  wire [15:0] _T_65206; // @[Mux.scala 19:72:@36853.4]
  wire [7:0] _T_65213; // @[Mux.scala 19:72:@36860.4]
  wire [7:0] _T_65220; // @[Mux.scala 19:72:@36867.4]
  wire [15:0] _T_65221; // @[Mux.scala 19:72:@36868.4]
  wire [15:0] _T_65223; // @[Mux.scala 19:72:@36869.4]
  wire [7:0] _T_65230; // @[Mux.scala 19:72:@36876.4]
  wire [7:0] _T_65237; // @[Mux.scala 19:72:@36883.4]
  wire [15:0] _T_65238; // @[Mux.scala 19:72:@36884.4]
  wire [15:0] _T_65240; // @[Mux.scala 19:72:@36885.4]
  wire [7:0] _T_65247; // @[Mux.scala 19:72:@36892.4]
  wire [7:0] _T_65254; // @[Mux.scala 19:72:@36899.4]
  wire [15:0] _T_65255; // @[Mux.scala 19:72:@36900.4]
  wire [15:0] _T_65257; // @[Mux.scala 19:72:@36901.4]
  wire [7:0] _T_65264; // @[Mux.scala 19:72:@36908.4]
  wire [7:0] _T_65271; // @[Mux.scala 19:72:@36915.4]
  wire [15:0] _T_65272; // @[Mux.scala 19:72:@36916.4]
  wire [15:0] _T_65274; // @[Mux.scala 19:72:@36917.4]
  wire [7:0] _T_65281; // @[Mux.scala 19:72:@36924.4]
  wire [7:0] _T_65288; // @[Mux.scala 19:72:@36931.4]
  wire [15:0] _T_65289; // @[Mux.scala 19:72:@36932.4]
  wire [15:0] _T_65291; // @[Mux.scala 19:72:@36933.4]
  wire [7:0] _T_65298; // @[Mux.scala 19:72:@36940.4]
  wire [7:0] _T_65305; // @[Mux.scala 19:72:@36947.4]
  wire [15:0] _T_65306; // @[Mux.scala 19:72:@36948.4]
  wire [15:0] _T_65308; // @[Mux.scala 19:72:@36949.4]
  wire [7:0] _T_65315; // @[Mux.scala 19:72:@36956.4]
  wire [7:0] _T_65322; // @[Mux.scala 19:72:@36963.4]
  wire [15:0] _T_65323; // @[Mux.scala 19:72:@36964.4]
  wire [15:0] _T_65325; // @[Mux.scala 19:72:@36965.4]
  wire [15:0] _T_65340; // @[Mux.scala 19:72:@36980.4]
  wire [15:0] _T_65342; // @[Mux.scala 19:72:@36981.4]
  wire [15:0] _T_65357; // @[Mux.scala 19:72:@36996.4]
  wire [15:0] _T_65359; // @[Mux.scala 19:72:@36997.4]
  wire [15:0] _T_65374; // @[Mux.scala 19:72:@37012.4]
  wire [15:0] _T_65376; // @[Mux.scala 19:72:@37013.4]
  wire [15:0] _T_65391; // @[Mux.scala 19:72:@37028.4]
  wire [15:0] _T_65393; // @[Mux.scala 19:72:@37029.4]
  wire [15:0] _T_65408; // @[Mux.scala 19:72:@37044.4]
  wire [15:0] _T_65410; // @[Mux.scala 19:72:@37045.4]
  wire [15:0] _T_65425; // @[Mux.scala 19:72:@37060.4]
  wire [15:0] _T_65427; // @[Mux.scala 19:72:@37061.4]
  wire [15:0] _T_65442; // @[Mux.scala 19:72:@37076.4]
  wire [15:0] _T_65444; // @[Mux.scala 19:72:@37077.4]
  wire [15:0] _T_65459; // @[Mux.scala 19:72:@37092.4]
  wire [15:0] _T_65461; // @[Mux.scala 19:72:@37093.4]
  wire [15:0] _T_65462; // @[Mux.scala 19:72:@37094.4]
  wire [15:0] _T_65463; // @[Mux.scala 19:72:@37095.4]
  wire [15:0] _T_65464; // @[Mux.scala 19:72:@37096.4]
  wire [15:0] _T_65465; // @[Mux.scala 19:72:@37097.4]
  wire [15:0] _T_65466; // @[Mux.scala 19:72:@37098.4]
  wire [15:0] _T_65467; // @[Mux.scala 19:72:@37099.4]
  wire [15:0] _T_65468; // @[Mux.scala 19:72:@37100.4]
  wire [15:0] _T_65469; // @[Mux.scala 19:72:@37101.4]
  wire [15:0] _T_65470; // @[Mux.scala 19:72:@37102.4]
  wire [15:0] _T_65471; // @[Mux.scala 19:72:@37103.4]
  wire [15:0] _T_65472; // @[Mux.scala 19:72:@37104.4]
  wire [15:0] _T_65473; // @[Mux.scala 19:72:@37105.4]
  wire [15:0] _T_65474; // @[Mux.scala 19:72:@37106.4]
  wire [15:0] _T_65475; // @[Mux.scala 19:72:@37107.4]
  wire [15:0] _T_65476; // @[Mux.scala 19:72:@37108.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_419;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_420;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_421;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_422;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_423;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_424;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_425;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_426;
  reg  storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_427;
  reg  storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_428;
  reg  storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_429;
  reg  storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_430;
  reg  storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_431;
  reg  storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_432;
  reg  storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_433;
  reg  storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_434;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_435;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_436;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_437;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_438;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_439;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_440;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_441;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_442;
  reg  storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_443;
  reg  storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_444;
  reg  storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_445;
  reg  storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_446;
  reg  storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_447;
  reg  storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_448;
  reg  storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_449;
  reg  storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_450;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_451;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_452;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_453;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_454;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_455;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_456;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_457;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_458;
  reg  storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_459;
  reg  storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_460;
  reg  storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_461;
  reg  storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_462;
  reg  storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_463;
  reg  storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_464;
  reg  storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_465;
  reg  storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_466;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_467;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_468;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_469;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_470;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_471;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_472;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_473;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_474;
  reg  storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_475;
  reg  storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_476;
  reg  storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_477;
  reg  storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_478;
  reg  storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_479;
  reg  storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_480;
  reg  storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_481;
  reg  storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_482;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_483;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_484;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_485;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_486;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_487;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_488;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_489;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_490;
  reg  storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_491;
  reg  storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_492;
  reg  storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_493;
  reg  storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_494;
  reg  storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_495;
  reg  storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_496;
  reg  storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_497;
  reg  storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_498;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_499;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_500;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_501;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_502;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_503;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_504;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_505;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_506;
  reg  storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_507;
  reg  storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_508;
  reg  storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_509;
  reg  storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_510;
  reg  storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_511;
  reg  storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_512;
  reg  storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_513;
  reg  storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_514;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_515;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_516;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_517;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_518;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_519;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_520;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_521;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_522;
  reg  storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_523;
  reg  storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_524;
  reg  storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_525;
  reg  storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_526;
  reg  storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_527;
  reg  storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_528;
  reg  storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_529;
  reg  storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_530;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_531;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_532;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_533;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_534;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_535;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_536;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_537;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_538;
  reg  storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_539;
  reg  storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_540;
  reg  storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_541;
  reg  storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_542;
  reg  storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_543;
  reg  storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_544;
  reg  storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_545;
  reg  storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_546;
  reg  storeAddrNotKnownFlagsPReg_8_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_547;
  reg  storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_548;
  reg  storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_549;
  reg  storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_550;
  reg  storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_551;
  reg  storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_552;
  reg  storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_553;
  reg  storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_554;
  reg  storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_555;
  reg  storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_556;
  reg  storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_557;
  reg  storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_558;
  reg  storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_559;
  reg  storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_560;
  reg  storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_561;
  reg  storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_562;
  reg  storeAddrNotKnownFlagsPReg_9_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_563;
  reg  storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_564;
  reg  storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_565;
  reg  storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_566;
  reg  storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_567;
  reg  storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_568;
  reg  storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_569;
  reg  storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_570;
  reg  storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_571;
  reg  storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_572;
  reg  storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_573;
  reg  storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_574;
  reg  storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_575;
  reg  storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_576;
  reg  storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_577;
  reg  storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_578;
  reg  storeAddrNotKnownFlagsPReg_10_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_579;
  reg  storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_580;
  reg  storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_581;
  reg  storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_582;
  reg  storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_583;
  reg  storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_584;
  reg  storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_585;
  reg  storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_586;
  reg  storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_587;
  reg  storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_588;
  reg  storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_589;
  reg  storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_590;
  reg  storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_591;
  reg  storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_592;
  reg  storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_593;
  reg  storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_594;
  reg  storeAddrNotKnownFlagsPReg_11_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_595;
  reg  storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_596;
  reg  storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_597;
  reg  storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_598;
  reg  storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_599;
  reg  storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_600;
  reg  storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_601;
  reg  storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_602;
  reg  storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_603;
  reg  storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_604;
  reg  storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_605;
  reg  storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_606;
  reg  storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_607;
  reg  storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_608;
  reg  storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_609;
  reg  storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_610;
  reg  storeAddrNotKnownFlagsPReg_12_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_611;
  reg  storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_612;
  reg  storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_613;
  reg  storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_614;
  reg  storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_615;
  reg  storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_616;
  reg  storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_617;
  reg  storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_618;
  reg  storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_619;
  reg  storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_620;
  reg  storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_621;
  reg  storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_622;
  reg  storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_623;
  reg  storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_624;
  reg  storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_625;
  reg  storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_626;
  reg  storeAddrNotKnownFlagsPReg_13_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_627;
  reg  storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_628;
  reg  storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_629;
  reg  storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_630;
  reg  storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_631;
  reg  storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_632;
  reg  storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_633;
  reg  storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_634;
  reg  storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_635;
  reg  storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_636;
  reg  storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_637;
  reg  storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_638;
  reg  storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_639;
  reg  storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_640;
  reg  storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_641;
  reg  storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_642;
  reg  storeAddrNotKnownFlagsPReg_14_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_643;
  reg  storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_644;
  reg  storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_645;
  reg  storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_646;
  reg  storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_647;
  reg  storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_648;
  reg  storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_649;
  reg  storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_650;
  reg  storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_651;
  reg  storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_652;
  reg  storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_653;
  reg  storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_654;
  reg  storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_655;
  reg  storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_656;
  reg  storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_657;
  reg  storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_658;
  reg  storeAddrNotKnownFlagsPReg_15_0; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_659;
  reg  storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_660;
  reg  storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_661;
  reg  storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_662;
  reg  storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_663;
  reg  storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_664;
  reg  storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_665;
  reg  storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_666;
  reg  storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_667;
  reg  storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_668;
  reg  storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_669;
  reg  storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_670;
  reg  storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_671;
  reg  storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_672;
  reg  storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_673;
  reg  storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 167:43:@37401.4]
  reg [31:0] _RAND_674;
  reg  shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_675;
  reg  shiftedStoreDataKnownPReg_1; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_676;
  reg  shiftedStoreDataKnownPReg_2; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_677;
  reg  shiftedStoreDataKnownPReg_3; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_678;
  reg  shiftedStoreDataKnownPReg_4; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_679;
  reg  shiftedStoreDataKnownPReg_5; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_680;
  reg  shiftedStoreDataKnownPReg_6; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_681;
  reg  shiftedStoreDataKnownPReg_7; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_682;
  reg  shiftedStoreDataKnownPReg_8; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_683;
  reg  shiftedStoreDataKnownPReg_9; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_684;
  reg  shiftedStoreDataKnownPReg_10; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_685;
  reg  shiftedStoreDataKnownPReg_11; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_686;
  reg  shiftedStoreDataKnownPReg_12; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_687;
  reg  shiftedStoreDataKnownPReg_13; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_688;
  reg  shiftedStoreDataKnownPReg_14; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_689;
  reg  shiftedStoreDataKnownPReg_15; // @[LoadQueue.scala 168:42:@37658.4]
  reg [31:0] _RAND_690;
  reg [31:0] shiftedStoreDataQPreg_0; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_691;
  reg [31:0] shiftedStoreDataQPreg_1; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_692;
  reg [31:0] shiftedStoreDataQPreg_2; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_693;
  reg [31:0] shiftedStoreDataQPreg_3; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_694;
  reg [31:0] shiftedStoreDataQPreg_4; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_695;
  reg [31:0] shiftedStoreDataQPreg_5; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_696;
  reg [31:0] shiftedStoreDataQPreg_6; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_697;
  reg [31:0] shiftedStoreDataQPreg_7; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_698;
  reg [31:0] shiftedStoreDataQPreg_8; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_699;
  reg [31:0] shiftedStoreDataQPreg_9; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_700;
  reg [31:0] shiftedStoreDataQPreg_10; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_701;
  reg [31:0] shiftedStoreDataQPreg_11; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_702;
  reg [31:0] shiftedStoreDataQPreg_12; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_703;
  reg [31:0] shiftedStoreDataQPreg_13; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_704;
  reg [31:0] shiftedStoreDataQPreg_14; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_705;
  reg [31:0] shiftedStoreDataQPreg_15; // @[LoadQueue.scala 169:38:@37675.4]
  reg [31:0] _RAND_706;
  reg  addrKnownPReg_0; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_707;
  reg  addrKnownPReg_1; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_708;
  reg  addrKnownPReg_2; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_709;
  reg  addrKnownPReg_3; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_710;
  reg  addrKnownPReg_4; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_711;
  reg  addrKnownPReg_5; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_712;
  reg  addrKnownPReg_6; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_713;
  reg  addrKnownPReg_7; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_714;
  reg  addrKnownPReg_8; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_715;
  reg  addrKnownPReg_9; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_716;
  reg  addrKnownPReg_10; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_717;
  reg  addrKnownPReg_11; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_718;
  reg  addrKnownPReg_12; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_719;
  reg  addrKnownPReg_13; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_720;
  reg  addrKnownPReg_14; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_721;
  reg  addrKnownPReg_15; // @[LoadQueue.scala 170:30:@37692.4]
  reg [31:0] _RAND_722;
  reg  dataKnownPReg_0; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_723;
  reg  dataKnownPReg_1; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_724;
  reg  dataKnownPReg_2; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_725;
  reg  dataKnownPReg_3; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_726;
  reg  dataKnownPReg_4; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_727;
  reg  dataKnownPReg_5; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_728;
  reg  dataKnownPReg_6; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_729;
  reg  dataKnownPReg_7; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_730;
  reg  dataKnownPReg_8; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_731;
  reg  dataKnownPReg_9; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_732;
  reg  dataKnownPReg_10; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_733;
  reg  dataKnownPReg_11; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_734;
  reg  dataKnownPReg_12; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_735;
  reg  dataKnownPReg_13; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_736;
  reg  dataKnownPReg_14; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_737;
  reg  dataKnownPReg_15; // @[LoadQueue.scala 171:30:@37709.4]
  reg [31:0] _RAND_738;
  wire [1:0] _T_88268; // @[LoadQueue.scala 191:60:@37781.4]
  wire [1:0] _T_88269; // @[LoadQueue.scala 191:60:@37782.4]
  wire [2:0] _T_88270; // @[LoadQueue.scala 191:60:@37783.4]
  wire [2:0] _T_88271; // @[LoadQueue.scala 191:60:@37784.4]
  wire [2:0] _T_88272; // @[LoadQueue.scala 191:60:@37785.4]
  wire [2:0] _T_88273; // @[LoadQueue.scala 191:60:@37786.4]
  wire [3:0] _T_88274; // @[LoadQueue.scala 191:60:@37787.4]
  wire [3:0] _T_88275; // @[LoadQueue.scala 191:60:@37788.4]
  wire [3:0] _T_88276; // @[LoadQueue.scala 191:60:@37789.4]
  wire [3:0] _T_88277; // @[LoadQueue.scala 191:60:@37790.4]
  wire [3:0] _T_88278; // @[LoadQueue.scala 191:60:@37791.4]
  wire [3:0] _T_88279; // @[LoadQueue.scala 191:60:@37792.4]
  wire [3:0] _T_88280; // @[LoadQueue.scala 191:60:@37793.4]
  wire [3:0] _T_88281; // @[LoadQueue.scala 191:60:@37794.4]
  wire  _T_88284; // @[LoadQueue.scala 192:43:@37796.4]
  wire  _T_88285; // @[LoadQueue.scala 192:43:@37797.4]
  wire  _T_88286; // @[LoadQueue.scala 192:43:@37798.4]
  wire  _T_88287; // @[LoadQueue.scala 192:43:@37799.4]
  wire  _T_88288; // @[LoadQueue.scala 192:43:@37800.4]
  wire  _T_88289; // @[LoadQueue.scala 192:43:@37801.4]
  wire  _T_88290; // @[LoadQueue.scala 192:43:@37802.4]
  wire  _T_88291; // @[LoadQueue.scala 192:43:@37803.4]
  wire  _T_88292; // @[LoadQueue.scala 192:43:@37804.4]
  wire  _T_88293; // @[LoadQueue.scala 192:43:@37805.4]
  wire  _T_88294; // @[LoadQueue.scala 192:43:@37806.4]
  wire  _T_88295; // @[LoadQueue.scala 192:43:@37807.4]
  wire  _T_88296; // @[LoadQueue.scala 192:43:@37808.4]
  wire  _T_88297; // @[LoadQueue.scala 192:43:@37809.4]
  wire  _T_88298; // @[LoadQueue.scala 192:43:@37810.4]
  wire  _GEN_864; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_865; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_866; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_867; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_868; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_869; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_870; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_871; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_872; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_873; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_874; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_875; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_876; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_877; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_878; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_879; // @[LoadQueue.scala 193:43:@37812.6]
  wire  _GEN_881; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_882; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_883; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_884; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_885; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_886; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_887; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_888; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_889; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_890; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_891; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_892; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_893; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_894; // @[LoadQueue.scala 194:31:@37813.6]
  wire  _GEN_895; // @[LoadQueue.scala 194:31:@37813.6]
  wire [31:0] _GEN_897; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_898; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_899; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_900; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_901; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_902; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_903; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_904; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_905; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_906; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_907; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_908; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_909; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_910; // @[LoadQueue.scala 195:31:@37814.6]
  wire [31:0] _GEN_911; // @[LoadQueue.scala 195:31:@37814.6]
  wire  lastConflict_0_0; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_1; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_2; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_3; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_4; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_5; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_6; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_7; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_8; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_9; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_10; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_11; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_12; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_13; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_14; // @[LoadQueue.scala 192:53:@37811.4]
  wire  lastConflict_0_15; // @[LoadQueue.scala 192:53:@37811.4]
  wire  canBypass_0; // @[LoadQueue.scala 192:53:@37811.4]
  wire [31:0] bypassVal_0; // @[LoadQueue.scala 192:53:@37811.4]
  wire [1:0] _T_88404; // @[LoadQueue.scala 191:60:@37868.4]
  wire [1:0] _T_88405; // @[LoadQueue.scala 191:60:@37869.4]
  wire [2:0] _T_88406; // @[LoadQueue.scala 191:60:@37870.4]
  wire [2:0] _T_88407; // @[LoadQueue.scala 191:60:@37871.4]
  wire [2:0] _T_88408; // @[LoadQueue.scala 191:60:@37872.4]
  wire [2:0] _T_88409; // @[LoadQueue.scala 191:60:@37873.4]
  wire [3:0] _T_88410; // @[LoadQueue.scala 191:60:@37874.4]
  wire [3:0] _T_88411; // @[LoadQueue.scala 191:60:@37875.4]
  wire [3:0] _T_88412; // @[LoadQueue.scala 191:60:@37876.4]
  wire [3:0] _T_88413; // @[LoadQueue.scala 191:60:@37877.4]
  wire [3:0] _T_88414; // @[LoadQueue.scala 191:60:@37878.4]
  wire [3:0] _T_88415; // @[LoadQueue.scala 191:60:@37879.4]
  wire [3:0] _T_88416; // @[LoadQueue.scala 191:60:@37880.4]
  wire [3:0] _T_88417; // @[LoadQueue.scala 191:60:@37881.4]
  wire  _T_88420; // @[LoadQueue.scala 192:43:@37883.4]
  wire  _T_88421; // @[LoadQueue.scala 192:43:@37884.4]
  wire  _T_88422; // @[LoadQueue.scala 192:43:@37885.4]
  wire  _T_88423; // @[LoadQueue.scala 192:43:@37886.4]
  wire  _T_88424; // @[LoadQueue.scala 192:43:@37887.4]
  wire  _T_88425; // @[LoadQueue.scala 192:43:@37888.4]
  wire  _T_88426; // @[LoadQueue.scala 192:43:@37889.4]
  wire  _T_88427; // @[LoadQueue.scala 192:43:@37890.4]
  wire  _T_88428; // @[LoadQueue.scala 192:43:@37891.4]
  wire  _T_88429; // @[LoadQueue.scala 192:43:@37892.4]
  wire  _T_88430; // @[LoadQueue.scala 192:43:@37893.4]
  wire  _T_88431; // @[LoadQueue.scala 192:43:@37894.4]
  wire  _T_88432; // @[LoadQueue.scala 192:43:@37895.4]
  wire  _T_88433; // @[LoadQueue.scala 192:43:@37896.4]
  wire  _T_88434; // @[LoadQueue.scala 192:43:@37897.4]
  wire  _GEN_930; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_931; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_932; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_933; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_934; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_935; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_936; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_937; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_938; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_939; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_940; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_941; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_942; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_943; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_944; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_945; // @[LoadQueue.scala 193:43:@37899.6]
  wire  _GEN_947; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_948; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_949; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_950; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_951; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_952; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_953; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_954; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_955; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_956; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_957; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_958; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_959; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_960; // @[LoadQueue.scala 194:31:@37900.6]
  wire  _GEN_961; // @[LoadQueue.scala 194:31:@37900.6]
  wire [31:0] _GEN_963; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_964; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_965; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_966; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_967; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_968; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_969; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_970; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_971; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_972; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_973; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_974; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_975; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_976; // @[LoadQueue.scala 195:31:@37901.6]
  wire [31:0] _GEN_977; // @[LoadQueue.scala 195:31:@37901.6]
  wire  lastConflict_1_0; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_1; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_2; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_3; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_4; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_5; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_6; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_7; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_8; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_9; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_10; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_11; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_12; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_13; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_14; // @[LoadQueue.scala 192:53:@37898.4]
  wire  lastConflict_1_15; // @[LoadQueue.scala 192:53:@37898.4]
  wire  canBypass_1; // @[LoadQueue.scala 192:53:@37898.4]
  wire [31:0] bypassVal_1; // @[LoadQueue.scala 192:53:@37898.4]
  wire [1:0] _T_88540; // @[LoadQueue.scala 191:60:@37955.4]
  wire [1:0] _T_88541; // @[LoadQueue.scala 191:60:@37956.4]
  wire [2:0] _T_88542; // @[LoadQueue.scala 191:60:@37957.4]
  wire [2:0] _T_88543; // @[LoadQueue.scala 191:60:@37958.4]
  wire [2:0] _T_88544; // @[LoadQueue.scala 191:60:@37959.4]
  wire [2:0] _T_88545; // @[LoadQueue.scala 191:60:@37960.4]
  wire [3:0] _T_88546; // @[LoadQueue.scala 191:60:@37961.4]
  wire [3:0] _T_88547; // @[LoadQueue.scala 191:60:@37962.4]
  wire [3:0] _T_88548; // @[LoadQueue.scala 191:60:@37963.4]
  wire [3:0] _T_88549; // @[LoadQueue.scala 191:60:@37964.4]
  wire [3:0] _T_88550; // @[LoadQueue.scala 191:60:@37965.4]
  wire [3:0] _T_88551; // @[LoadQueue.scala 191:60:@37966.4]
  wire [3:0] _T_88552; // @[LoadQueue.scala 191:60:@37967.4]
  wire [3:0] _T_88553; // @[LoadQueue.scala 191:60:@37968.4]
  wire  _T_88556; // @[LoadQueue.scala 192:43:@37970.4]
  wire  _T_88557; // @[LoadQueue.scala 192:43:@37971.4]
  wire  _T_88558; // @[LoadQueue.scala 192:43:@37972.4]
  wire  _T_88559; // @[LoadQueue.scala 192:43:@37973.4]
  wire  _T_88560; // @[LoadQueue.scala 192:43:@37974.4]
  wire  _T_88561; // @[LoadQueue.scala 192:43:@37975.4]
  wire  _T_88562; // @[LoadQueue.scala 192:43:@37976.4]
  wire  _T_88563; // @[LoadQueue.scala 192:43:@37977.4]
  wire  _T_88564; // @[LoadQueue.scala 192:43:@37978.4]
  wire  _T_88565; // @[LoadQueue.scala 192:43:@37979.4]
  wire  _T_88566; // @[LoadQueue.scala 192:43:@37980.4]
  wire  _T_88567; // @[LoadQueue.scala 192:43:@37981.4]
  wire  _T_88568; // @[LoadQueue.scala 192:43:@37982.4]
  wire  _T_88569; // @[LoadQueue.scala 192:43:@37983.4]
  wire  _T_88570; // @[LoadQueue.scala 192:43:@37984.4]
  wire  _GEN_996; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_997; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_998; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_999; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1000; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1001; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1002; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1003; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1004; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1005; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1006; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1007; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1008; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1009; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1010; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1011; // @[LoadQueue.scala 193:43:@37986.6]
  wire  _GEN_1013; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1014; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1015; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1016; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1017; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1018; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1019; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1020; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1021; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1022; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1023; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1024; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1025; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1026; // @[LoadQueue.scala 194:31:@37987.6]
  wire  _GEN_1027; // @[LoadQueue.scala 194:31:@37987.6]
  wire [31:0] _GEN_1029; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1030; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1031; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1032; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1033; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1034; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1035; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1036; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1037; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1038; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1039; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1040; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1041; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1042; // @[LoadQueue.scala 195:31:@37988.6]
  wire [31:0] _GEN_1043; // @[LoadQueue.scala 195:31:@37988.6]
  wire  lastConflict_2_0; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_1; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_2; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_3; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_4; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_5; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_6; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_7; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_8; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_9; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_10; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_11; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_12; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_13; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_14; // @[LoadQueue.scala 192:53:@37985.4]
  wire  lastConflict_2_15; // @[LoadQueue.scala 192:53:@37985.4]
  wire  canBypass_2; // @[LoadQueue.scala 192:53:@37985.4]
  wire [31:0] bypassVal_2; // @[LoadQueue.scala 192:53:@37985.4]
  wire [1:0] _T_88676; // @[LoadQueue.scala 191:60:@38042.4]
  wire [1:0] _T_88677; // @[LoadQueue.scala 191:60:@38043.4]
  wire [2:0] _T_88678; // @[LoadQueue.scala 191:60:@38044.4]
  wire [2:0] _T_88679; // @[LoadQueue.scala 191:60:@38045.4]
  wire [2:0] _T_88680; // @[LoadQueue.scala 191:60:@38046.4]
  wire [2:0] _T_88681; // @[LoadQueue.scala 191:60:@38047.4]
  wire [3:0] _T_88682; // @[LoadQueue.scala 191:60:@38048.4]
  wire [3:0] _T_88683; // @[LoadQueue.scala 191:60:@38049.4]
  wire [3:0] _T_88684; // @[LoadQueue.scala 191:60:@38050.4]
  wire [3:0] _T_88685; // @[LoadQueue.scala 191:60:@38051.4]
  wire [3:0] _T_88686; // @[LoadQueue.scala 191:60:@38052.4]
  wire [3:0] _T_88687; // @[LoadQueue.scala 191:60:@38053.4]
  wire [3:0] _T_88688; // @[LoadQueue.scala 191:60:@38054.4]
  wire [3:0] _T_88689; // @[LoadQueue.scala 191:60:@38055.4]
  wire  _T_88692; // @[LoadQueue.scala 192:43:@38057.4]
  wire  _T_88693; // @[LoadQueue.scala 192:43:@38058.4]
  wire  _T_88694; // @[LoadQueue.scala 192:43:@38059.4]
  wire  _T_88695; // @[LoadQueue.scala 192:43:@38060.4]
  wire  _T_88696; // @[LoadQueue.scala 192:43:@38061.4]
  wire  _T_88697; // @[LoadQueue.scala 192:43:@38062.4]
  wire  _T_88698; // @[LoadQueue.scala 192:43:@38063.4]
  wire  _T_88699; // @[LoadQueue.scala 192:43:@38064.4]
  wire  _T_88700; // @[LoadQueue.scala 192:43:@38065.4]
  wire  _T_88701; // @[LoadQueue.scala 192:43:@38066.4]
  wire  _T_88702; // @[LoadQueue.scala 192:43:@38067.4]
  wire  _T_88703; // @[LoadQueue.scala 192:43:@38068.4]
  wire  _T_88704; // @[LoadQueue.scala 192:43:@38069.4]
  wire  _T_88705; // @[LoadQueue.scala 192:43:@38070.4]
  wire  _T_88706; // @[LoadQueue.scala 192:43:@38071.4]
  wire  _GEN_1062; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1063; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1064; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1065; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1066; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1067; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1068; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1069; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1070; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1071; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1072; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1073; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1074; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1075; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1076; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1077; // @[LoadQueue.scala 193:43:@38073.6]
  wire  _GEN_1079; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1080; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1081; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1082; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1083; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1084; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1085; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1086; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1087; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1088; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1089; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1090; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1091; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1092; // @[LoadQueue.scala 194:31:@38074.6]
  wire  _GEN_1093; // @[LoadQueue.scala 194:31:@38074.6]
  wire [31:0] _GEN_1095; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1096; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1097; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1098; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1099; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1100; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1101; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1102; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1103; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1104; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1105; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1106; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1107; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1108; // @[LoadQueue.scala 195:31:@38075.6]
  wire [31:0] _GEN_1109; // @[LoadQueue.scala 195:31:@38075.6]
  wire  lastConflict_3_0; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_1; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_2; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_3; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_4; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_5; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_6; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_7; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_8; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_9; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_10; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_11; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_12; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_13; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_14; // @[LoadQueue.scala 192:53:@38072.4]
  wire  lastConflict_3_15; // @[LoadQueue.scala 192:53:@38072.4]
  wire  canBypass_3; // @[LoadQueue.scala 192:53:@38072.4]
  wire [31:0] bypassVal_3; // @[LoadQueue.scala 192:53:@38072.4]
  wire [1:0] _T_88812; // @[LoadQueue.scala 191:60:@38129.4]
  wire [1:0] _T_88813; // @[LoadQueue.scala 191:60:@38130.4]
  wire [2:0] _T_88814; // @[LoadQueue.scala 191:60:@38131.4]
  wire [2:0] _T_88815; // @[LoadQueue.scala 191:60:@38132.4]
  wire [2:0] _T_88816; // @[LoadQueue.scala 191:60:@38133.4]
  wire [2:0] _T_88817; // @[LoadQueue.scala 191:60:@38134.4]
  wire [3:0] _T_88818; // @[LoadQueue.scala 191:60:@38135.4]
  wire [3:0] _T_88819; // @[LoadQueue.scala 191:60:@38136.4]
  wire [3:0] _T_88820; // @[LoadQueue.scala 191:60:@38137.4]
  wire [3:0] _T_88821; // @[LoadQueue.scala 191:60:@38138.4]
  wire [3:0] _T_88822; // @[LoadQueue.scala 191:60:@38139.4]
  wire [3:0] _T_88823; // @[LoadQueue.scala 191:60:@38140.4]
  wire [3:0] _T_88824; // @[LoadQueue.scala 191:60:@38141.4]
  wire [3:0] _T_88825; // @[LoadQueue.scala 191:60:@38142.4]
  wire  _T_88828; // @[LoadQueue.scala 192:43:@38144.4]
  wire  _T_88829; // @[LoadQueue.scala 192:43:@38145.4]
  wire  _T_88830; // @[LoadQueue.scala 192:43:@38146.4]
  wire  _T_88831; // @[LoadQueue.scala 192:43:@38147.4]
  wire  _T_88832; // @[LoadQueue.scala 192:43:@38148.4]
  wire  _T_88833; // @[LoadQueue.scala 192:43:@38149.4]
  wire  _T_88834; // @[LoadQueue.scala 192:43:@38150.4]
  wire  _T_88835; // @[LoadQueue.scala 192:43:@38151.4]
  wire  _T_88836; // @[LoadQueue.scala 192:43:@38152.4]
  wire  _T_88837; // @[LoadQueue.scala 192:43:@38153.4]
  wire  _T_88838; // @[LoadQueue.scala 192:43:@38154.4]
  wire  _T_88839; // @[LoadQueue.scala 192:43:@38155.4]
  wire  _T_88840; // @[LoadQueue.scala 192:43:@38156.4]
  wire  _T_88841; // @[LoadQueue.scala 192:43:@38157.4]
  wire  _T_88842; // @[LoadQueue.scala 192:43:@38158.4]
  wire  _GEN_1128; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1129; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1130; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1131; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1132; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1133; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1134; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1135; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1136; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1137; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1138; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1139; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1140; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1141; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1142; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1143; // @[LoadQueue.scala 193:43:@38160.6]
  wire  _GEN_1145; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1146; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1147; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1148; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1149; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1150; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1151; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1152; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1153; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1154; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1155; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1156; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1157; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1158; // @[LoadQueue.scala 194:31:@38161.6]
  wire  _GEN_1159; // @[LoadQueue.scala 194:31:@38161.6]
  wire [31:0] _GEN_1161; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1162; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1163; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1164; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1165; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1166; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1167; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1168; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1169; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1170; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1171; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1172; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1173; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1174; // @[LoadQueue.scala 195:31:@38162.6]
  wire [31:0] _GEN_1175; // @[LoadQueue.scala 195:31:@38162.6]
  wire  lastConflict_4_0; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_1; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_2; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_3; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_4; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_5; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_6; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_7; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_8; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_9; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_10; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_11; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_12; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_13; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_14; // @[LoadQueue.scala 192:53:@38159.4]
  wire  lastConflict_4_15; // @[LoadQueue.scala 192:53:@38159.4]
  wire  canBypass_4; // @[LoadQueue.scala 192:53:@38159.4]
  wire [31:0] bypassVal_4; // @[LoadQueue.scala 192:53:@38159.4]
  wire [1:0] _T_88948; // @[LoadQueue.scala 191:60:@38216.4]
  wire [1:0] _T_88949; // @[LoadQueue.scala 191:60:@38217.4]
  wire [2:0] _T_88950; // @[LoadQueue.scala 191:60:@38218.4]
  wire [2:0] _T_88951; // @[LoadQueue.scala 191:60:@38219.4]
  wire [2:0] _T_88952; // @[LoadQueue.scala 191:60:@38220.4]
  wire [2:0] _T_88953; // @[LoadQueue.scala 191:60:@38221.4]
  wire [3:0] _T_88954; // @[LoadQueue.scala 191:60:@38222.4]
  wire [3:0] _T_88955; // @[LoadQueue.scala 191:60:@38223.4]
  wire [3:0] _T_88956; // @[LoadQueue.scala 191:60:@38224.4]
  wire [3:0] _T_88957; // @[LoadQueue.scala 191:60:@38225.4]
  wire [3:0] _T_88958; // @[LoadQueue.scala 191:60:@38226.4]
  wire [3:0] _T_88959; // @[LoadQueue.scala 191:60:@38227.4]
  wire [3:0] _T_88960; // @[LoadQueue.scala 191:60:@38228.4]
  wire [3:0] _T_88961; // @[LoadQueue.scala 191:60:@38229.4]
  wire  _T_88964; // @[LoadQueue.scala 192:43:@38231.4]
  wire  _T_88965; // @[LoadQueue.scala 192:43:@38232.4]
  wire  _T_88966; // @[LoadQueue.scala 192:43:@38233.4]
  wire  _T_88967; // @[LoadQueue.scala 192:43:@38234.4]
  wire  _T_88968; // @[LoadQueue.scala 192:43:@38235.4]
  wire  _T_88969; // @[LoadQueue.scala 192:43:@38236.4]
  wire  _T_88970; // @[LoadQueue.scala 192:43:@38237.4]
  wire  _T_88971; // @[LoadQueue.scala 192:43:@38238.4]
  wire  _T_88972; // @[LoadQueue.scala 192:43:@38239.4]
  wire  _T_88973; // @[LoadQueue.scala 192:43:@38240.4]
  wire  _T_88974; // @[LoadQueue.scala 192:43:@38241.4]
  wire  _T_88975; // @[LoadQueue.scala 192:43:@38242.4]
  wire  _T_88976; // @[LoadQueue.scala 192:43:@38243.4]
  wire  _T_88977; // @[LoadQueue.scala 192:43:@38244.4]
  wire  _T_88978; // @[LoadQueue.scala 192:43:@38245.4]
  wire  _GEN_1194; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1195; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1196; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1197; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1198; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1199; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1200; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1201; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1202; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1203; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1204; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1205; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1206; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1207; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1208; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1209; // @[LoadQueue.scala 193:43:@38247.6]
  wire  _GEN_1211; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1212; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1213; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1214; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1215; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1216; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1217; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1218; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1219; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1220; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1221; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1222; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1223; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1224; // @[LoadQueue.scala 194:31:@38248.6]
  wire  _GEN_1225; // @[LoadQueue.scala 194:31:@38248.6]
  wire [31:0] _GEN_1227; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1228; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1229; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1230; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1231; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1232; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1233; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1234; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1235; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1236; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1237; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1238; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1239; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1240; // @[LoadQueue.scala 195:31:@38249.6]
  wire [31:0] _GEN_1241; // @[LoadQueue.scala 195:31:@38249.6]
  wire  lastConflict_5_0; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_1; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_2; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_3; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_4; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_5; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_6; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_7; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_8; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_9; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_10; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_11; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_12; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_13; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_14; // @[LoadQueue.scala 192:53:@38246.4]
  wire  lastConflict_5_15; // @[LoadQueue.scala 192:53:@38246.4]
  wire  canBypass_5; // @[LoadQueue.scala 192:53:@38246.4]
  wire [31:0] bypassVal_5; // @[LoadQueue.scala 192:53:@38246.4]
  wire [1:0] _T_89084; // @[LoadQueue.scala 191:60:@38303.4]
  wire [1:0] _T_89085; // @[LoadQueue.scala 191:60:@38304.4]
  wire [2:0] _T_89086; // @[LoadQueue.scala 191:60:@38305.4]
  wire [2:0] _T_89087; // @[LoadQueue.scala 191:60:@38306.4]
  wire [2:0] _T_89088; // @[LoadQueue.scala 191:60:@38307.4]
  wire [2:0] _T_89089; // @[LoadQueue.scala 191:60:@38308.4]
  wire [3:0] _T_89090; // @[LoadQueue.scala 191:60:@38309.4]
  wire [3:0] _T_89091; // @[LoadQueue.scala 191:60:@38310.4]
  wire [3:0] _T_89092; // @[LoadQueue.scala 191:60:@38311.4]
  wire [3:0] _T_89093; // @[LoadQueue.scala 191:60:@38312.4]
  wire [3:0] _T_89094; // @[LoadQueue.scala 191:60:@38313.4]
  wire [3:0] _T_89095; // @[LoadQueue.scala 191:60:@38314.4]
  wire [3:0] _T_89096; // @[LoadQueue.scala 191:60:@38315.4]
  wire [3:0] _T_89097; // @[LoadQueue.scala 191:60:@38316.4]
  wire  _T_89100; // @[LoadQueue.scala 192:43:@38318.4]
  wire  _T_89101; // @[LoadQueue.scala 192:43:@38319.4]
  wire  _T_89102; // @[LoadQueue.scala 192:43:@38320.4]
  wire  _T_89103; // @[LoadQueue.scala 192:43:@38321.4]
  wire  _T_89104; // @[LoadQueue.scala 192:43:@38322.4]
  wire  _T_89105; // @[LoadQueue.scala 192:43:@38323.4]
  wire  _T_89106; // @[LoadQueue.scala 192:43:@38324.4]
  wire  _T_89107; // @[LoadQueue.scala 192:43:@38325.4]
  wire  _T_89108; // @[LoadQueue.scala 192:43:@38326.4]
  wire  _T_89109; // @[LoadQueue.scala 192:43:@38327.4]
  wire  _T_89110; // @[LoadQueue.scala 192:43:@38328.4]
  wire  _T_89111; // @[LoadQueue.scala 192:43:@38329.4]
  wire  _T_89112; // @[LoadQueue.scala 192:43:@38330.4]
  wire  _T_89113; // @[LoadQueue.scala 192:43:@38331.4]
  wire  _T_89114; // @[LoadQueue.scala 192:43:@38332.4]
  wire  _GEN_1260; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1261; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1262; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1263; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1264; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1265; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1266; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1267; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1268; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1269; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1270; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1271; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1272; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1273; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1274; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1275; // @[LoadQueue.scala 193:43:@38334.6]
  wire  _GEN_1277; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1278; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1279; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1280; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1281; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1282; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1283; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1284; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1285; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1286; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1287; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1288; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1289; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1290; // @[LoadQueue.scala 194:31:@38335.6]
  wire  _GEN_1291; // @[LoadQueue.scala 194:31:@38335.6]
  wire [31:0] _GEN_1293; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1294; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1295; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1296; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1297; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1298; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1299; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1300; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1301; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1302; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1303; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1304; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1305; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1306; // @[LoadQueue.scala 195:31:@38336.6]
  wire [31:0] _GEN_1307; // @[LoadQueue.scala 195:31:@38336.6]
  wire  lastConflict_6_0; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_1; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_2; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_3; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_4; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_5; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_6; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_7; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_8; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_9; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_10; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_11; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_12; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_13; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_14; // @[LoadQueue.scala 192:53:@38333.4]
  wire  lastConflict_6_15; // @[LoadQueue.scala 192:53:@38333.4]
  wire  canBypass_6; // @[LoadQueue.scala 192:53:@38333.4]
  wire [31:0] bypassVal_6; // @[LoadQueue.scala 192:53:@38333.4]
  wire [1:0] _T_89220; // @[LoadQueue.scala 191:60:@38390.4]
  wire [1:0] _T_89221; // @[LoadQueue.scala 191:60:@38391.4]
  wire [2:0] _T_89222; // @[LoadQueue.scala 191:60:@38392.4]
  wire [2:0] _T_89223; // @[LoadQueue.scala 191:60:@38393.4]
  wire [2:0] _T_89224; // @[LoadQueue.scala 191:60:@38394.4]
  wire [2:0] _T_89225; // @[LoadQueue.scala 191:60:@38395.4]
  wire [3:0] _T_89226; // @[LoadQueue.scala 191:60:@38396.4]
  wire [3:0] _T_89227; // @[LoadQueue.scala 191:60:@38397.4]
  wire [3:0] _T_89228; // @[LoadQueue.scala 191:60:@38398.4]
  wire [3:0] _T_89229; // @[LoadQueue.scala 191:60:@38399.4]
  wire [3:0] _T_89230; // @[LoadQueue.scala 191:60:@38400.4]
  wire [3:0] _T_89231; // @[LoadQueue.scala 191:60:@38401.4]
  wire [3:0] _T_89232; // @[LoadQueue.scala 191:60:@38402.4]
  wire [3:0] _T_89233; // @[LoadQueue.scala 191:60:@38403.4]
  wire  _T_89236; // @[LoadQueue.scala 192:43:@38405.4]
  wire  _T_89237; // @[LoadQueue.scala 192:43:@38406.4]
  wire  _T_89238; // @[LoadQueue.scala 192:43:@38407.4]
  wire  _T_89239; // @[LoadQueue.scala 192:43:@38408.4]
  wire  _T_89240; // @[LoadQueue.scala 192:43:@38409.4]
  wire  _T_89241; // @[LoadQueue.scala 192:43:@38410.4]
  wire  _T_89242; // @[LoadQueue.scala 192:43:@38411.4]
  wire  _T_89243; // @[LoadQueue.scala 192:43:@38412.4]
  wire  _T_89244; // @[LoadQueue.scala 192:43:@38413.4]
  wire  _T_89245; // @[LoadQueue.scala 192:43:@38414.4]
  wire  _T_89246; // @[LoadQueue.scala 192:43:@38415.4]
  wire  _T_89247; // @[LoadQueue.scala 192:43:@38416.4]
  wire  _T_89248; // @[LoadQueue.scala 192:43:@38417.4]
  wire  _T_89249; // @[LoadQueue.scala 192:43:@38418.4]
  wire  _T_89250; // @[LoadQueue.scala 192:43:@38419.4]
  wire  _GEN_1326; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1327; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1328; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1329; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1330; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1331; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1332; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1333; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1334; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1335; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1336; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1337; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1338; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1339; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1340; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1341; // @[LoadQueue.scala 193:43:@38421.6]
  wire  _GEN_1343; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1344; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1345; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1346; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1347; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1348; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1349; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1350; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1351; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1352; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1353; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1354; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1355; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1356; // @[LoadQueue.scala 194:31:@38422.6]
  wire  _GEN_1357; // @[LoadQueue.scala 194:31:@38422.6]
  wire [31:0] _GEN_1359; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1360; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1361; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1362; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1363; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1364; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1365; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1366; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1367; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1368; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1369; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1370; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1371; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1372; // @[LoadQueue.scala 195:31:@38423.6]
  wire [31:0] _GEN_1373; // @[LoadQueue.scala 195:31:@38423.6]
  wire  lastConflict_7_0; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_1; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_2; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_3; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_4; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_5; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_6; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_7; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_8; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_9; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_10; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_11; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_12; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_13; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_14; // @[LoadQueue.scala 192:53:@38420.4]
  wire  lastConflict_7_15; // @[LoadQueue.scala 192:53:@38420.4]
  wire  canBypass_7; // @[LoadQueue.scala 192:53:@38420.4]
  wire [31:0] bypassVal_7; // @[LoadQueue.scala 192:53:@38420.4]
  wire [1:0] _T_89356; // @[LoadQueue.scala 191:60:@38477.4]
  wire [1:0] _T_89357; // @[LoadQueue.scala 191:60:@38478.4]
  wire [2:0] _T_89358; // @[LoadQueue.scala 191:60:@38479.4]
  wire [2:0] _T_89359; // @[LoadQueue.scala 191:60:@38480.4]
  wire [2:0] _T_89360; // @[LoadQueue.scala 191:60:@38481.4]
  wire [2:0] _T_89361; // @[LoadQueue.scala 191:60:@38482.4]
  wire [3:0] _T_89362; // @[LoadQueue.scala 191:60:@38483.4]
  wire [3:0] _T_89363; // @[LoadQueue.scala 191:60:@38484.4]
  wire [3:0] _T_89364; // @[LoadQueue.scala 191:60:@38485.4]
  wire [3:0] _T_89365; // @[LoadQueue.scala 191:60:@38486.4]
  wire [3:0] _T_89366; // @[LoadQueue.scala 191:60:@38487.4]
  wire [3:0] _T_89367; // @[LoadQueue.scala 191:60:@38488.4]
  wire [3:0] _T_89368; // @[LoadQueue.scala 191:60:@38489.4]
  wire [3:0] _T_89369; // @[LoadQueue.scala 191:60:@38490.4]
  wire  _T_89372; // @[LoadQueue.scala 192:43:@38492.4]
  wire  _T_89373; // @[LoadQueue.scala 192:43:@38493.4]
  wire  _T_89374; // @[LoadQueue.scala 192:43:@38494.4]
  wire  _T_89375; // @[LoadQueue.scala 192:43:@38495.4]
  wire  _T_89376; // @[LoadQueue.scala 192:43:@38496.4]
  wire  _T_89377; // @[LoadQueue.scala 192:43:@38497.4]
  wire  _T_89378; // @[LoadQueue.scala 192:43:@38498.4]
  wire  _T_89379; // @[LoadQueue.scala 192:43:@38499.4]
  wire  _T_89380; // @[LoadQueue.scala 192:43:@38500.4]
  wire  _T_89381; // @[LoadQueue.scala 192:43:@38501.4]
  wire  _T_89382; // @[LoadQueue.scala 192:43:@38502.4]
  wire  _T_89383; // @[LoadQueue.scala 192:43:@38503.4]
  wire  _T_89384; // @[LoadQueue.scala 192:43:@38504.4]
  wire  _T_89385; // @[LoadQueue.scala 192:43:@38505.4]
  wire  _T_89386; // @[LoadQueue.scala 192:43:@38506.4]
  wire  _GEN_1392; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1393; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1394; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1395; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1396; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1397; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1398; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1399; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1400; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1401; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1402; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1403; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1404; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1405; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1406; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1407; // @[LoadQueue.scala 193:43:@38508.6]
  wire  _GEN_1409; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1410; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1411; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1412; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1413; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1414; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1415; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1416; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1417; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1418; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1419; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1420; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1421; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1422; // @[LoadQueue.scala 194:31:@38509.6]
  wire  _GEN_1423; // @[LoadQueue.scala 194:31:@38509.6]
  wire [31:0] _GEN_1425; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1426; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1427; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1428; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1429; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1430; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1431; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1432; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1433; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1434; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1435; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1436; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1437; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1438; // @[LoadQueue.scala 195:31:@38510.6]
  wire [31:0] _GEN_1439; // @[LoadQueue.scala 195:31:@38510.6]
  wire  lastConflict_8_0; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_1; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_2; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_3; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_4; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_5; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_6; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_7; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_8; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_9; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_10; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_11; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_12; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_13; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_14; // @[LoadQueue.scala 192:53:@38507.4]
  wire  lastConflict_8_15; // @[LoadQueue.scala 192:53:@38507.4]
  wire  canBypass_8; // @[LoadQueue.scala 192:53:@38507.4]
  wire [31:0] bypassVal_8; // @[LoadQueue.scala 192:53:@38507.4]
  wire [1:0] _T_89492; // @[LoadQueue.scala 191:60:@38564.4]
  wire [1:0] _T_89493; // @[LoadQueue.scala 191:60:@38565.4]
  wire [2:0] _T_89494; // @[LoadQueue.scala 191:60:@38566.4]
  wire [2:0] _T_89495; // @[LoadQueue.scala 191:60:@38567.4]
  wire [2:0] _T_89496; // @[LoadQueue.scala 191:60:@38568.4]
  wire [2:0] _T_89497; // @[LoadQueue.scala 191:60:@38569.4]
  wire [3:0] _T_89498; // @[LoadQueue.scala 191:60:@38570.4]
  wire [3:0] _T_89499; // @[LoadQueue.scala 191:60:@38571.4]
  wire [3:0] _T_89500; // @[LoadQueue.scala 191:60:@38572.4]
  wire [3:0] _T_89501; // @[LoadQueue.scala 191:60:@38573.4]
  wire [3:0] _T_89502; // @[LoadQueue.scala 191:60:@38574.4]
  wire [3:0] _T_89503; // @[LoadQueue.scala 191:60:@38575.4]
  wire [3:0] _T_89504; // @[LoadQueue.scala 191:60:@38576.4]
  wire [3:0] _T_89505; // @[LoadQueue.scala 191:60:@38577.4]
  wire  _T_89508; // @[LoadQueue.scala 192:43:@38579.4]
  wire  _T_89509; // @[LoadQueue.scala 192:43:@38580.4]
  wire  _T_89510; // @[LoadQueue.scala 192:43:@38581.4]
  wire  _T_89511; // @[LoadQueue.scala 192:43:@38582.4]
  wire  _T_89512; // @[LoadQueue.scala 192:43:@38583.4]
  wire  _T_89513; // @[LoadQueue.scala 192:43:@38584.4]
  wire  _T_89514; // @[LoadQueue.scala 192:43:@38585.4]
  wire  _T_89515; // @[LoadQueue.scala 192:43:@38586.4]
  wire  _T_89516; // @[LoadQueue.scala 192:43:@38587.4]
  wire  _T_89517; // @[LoadQueue.scala 192:43:@38588.4]
  wire  _T_89518; // @[LoadQueue.scala 192:43:@38589.4]
  wire  _T_89519; // @[LoadQueue.scala 192:43:@38590.4]
  wire  _T_89520; // @[LoadQueue.scala 192:43:@38591.4]
  wire  _T_89521; // @[LoadQueue.scala 192:43:@38592.4]
  wire  _T_89522; // @[LoadQueue.scala 192:43:@38593.4]
  wire  _GEN_1458; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1459; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1460; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1461; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1462; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1463; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1464; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1465; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1466; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1467; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1468; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1469; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1470; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1471; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1472; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1473; // @[LoadQueue.scala 193:43:@38595.6]
  wire  _GEN_1475; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1476; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1477; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1478; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1479; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1480; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1481; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1482; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1483; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1484; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1485; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1486; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1487; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1488; // @[LoadQueue.scala 194:31:@38596.6]
  wire  _GEN_1489; // @[LoadQueue.scala 194:31:@38596.6]
  wire [31:0] _GEN_1491; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1492; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1493; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1494; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1495; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1496; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1497; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1498; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1499; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1500; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1501; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1502; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1503; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1504; // @[LoadQueue.scala 195:31:@38597.6]
  wire [31:0] _GEN_1505; // @[LoadQueue.scala 195:31:@38597.6]
  wire  lastConflict_9_0; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_1; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_2; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_3; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_4; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_5; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_6; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_7; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_8; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_9; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_10; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_11; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_12; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_13; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_14; // @[LoadQueue.scala 192:53:@38594.4]
  wire  lastConflict_9_15; // @[LoadQueue.scala 192:53:@38594.4]
  wire  canBypass_9; // @[LoadQueue.scala 192:53:@38594.4]
  wire [31:0] bypassVal_9; // @[LoadQueue.scala 192:53:@38594.4]
  wire [1:0] _T_89628; // @[LoadQueue.scala 191:60:@38651.4]
  wire [1:0] _T_89629; // @[LoadQueue.scala 191:60:@38652.4]
  wire [2:0] _T_89630; // @[LoadQueue.scala 191:60:@38653.4]
  wire [2:0] _T_89631; // @[LoadQueue.scala 191:60:@38654.4]
  wire [2:0] _T_89632; // @[LoadQueue.scala 191:60:@38655.4]
  wire [2:0] _T_89633; // @[LoadQueue.scala 191:60:@38656.4]
  wire [3:0] _T_89634; // @[LoadQueue.scala 191:60:@38657.4]
  wire [3:0] _T_89635; // @[LoadQueue.scala 191:60:@38658.4]
  wire [3:0] _T_89636; // @[LoadQueue.scala 191:60:@38659.4]
  wire [3:0] _T_89637; // @[LoadQueue.scala 191:60:@38660.4]
  wire [3:0] _T_89638; // @[LoadQueue.scala 191:60:@38661.4]
  wire [3:0] _T_89639; // @[LoadQueue.scala 191:60:@38662.4]
  wire [3:0] _T_89640; // @[LoadQueue.scala 191:60:@38663.4]
  wire [3:0] _T_89641; // @[LoadQueue.scala 191:60:@38664.4]
  wire  _T_89644; // @[LoadQueue.scala 192:43:@38666.4]
  wire  _T_89645; // @[LoadQueue.scala 192:43:@38667.4]
  wire  _T_89646; // @[LoadQueue.scala 192:43:@38668.4]
  wire  _T_89647; // @[LoadQueue.scala 192:43:@38669.4]
  wire  _T_89648; // @[LoadQueue.scala 192:43:@38670.4]
  wire  _T_89649; // @[LoadQueue.scala 192:43:@38671.4]
  wire  _T_89650; // @[LoadQueue.scala 192:43:@38672.4]
  wire  _T_89651; // @[LoadQueue.scala 192:43:@38673.4]
  wire  _T_89652; // @[LoadQueue.scala 192:43:@38674.4]
  wire  _T_89653; // @[LoadQueue.scala 192:43:@38675.4]
  wire  _T_89654; // @[LoadQueue.scala 192:43:@38676.4]
  wire  _T_89655; // @[LoadQueue.scala 192:43:@38677.4]
  wire  _T_89656; // @[LoadQueue.scala 192:43:@38678.4]
  wire  _T_89657; // @[LoadQueue.scala 192:43:@38679.4]
  wire  _T_89658; // @[LoadQueue.scala 192:43:@38680.4]
  wire  _GEN_1524; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1525; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1526; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1527; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1528; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1529; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1530; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1531; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1532; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1533; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1534; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1535; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1536; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1537; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1538; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1539; // @[LoadQueue.scala 193:43:@38682.6]
  wire  _GEN_1541; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1542; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1543; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1544; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1545; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1546; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1547; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1548; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1549; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1550; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1551; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1552; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1553; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1554; // @[LoadQueue.scala 194:31:@38683.6]
  wire  _GEN_1555; // @[LoadQueue.scala 194:31:@38683.6]
  wire [31:0] _GEN_1557; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1558; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1559; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1560; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1561; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1562; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1563; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1564; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1565; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1566; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1567; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1568; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1569; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1570; // @[LoadQueue.scala 195:31:@38684.6]
  wire [31:0] _GEN_1571; // @[LoadQueue.scala 195:31:@38684.6]
  wire  lastConflict_10_0; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_1; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_2; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_3; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_4; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_5; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_6; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_7; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_8; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_9; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_10; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_11; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_12; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_13; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_14; // @[LoadQueue.scala 192:53:@38681.4]
  wire  lastConflict_10_15; // @[LoadQueue.scala 192:53:@38681.4]
  wire  canBypass_10; // @[LoadQueue.scala 192:53:@38681.4]
  wire [31:0] bypassVal_10; // @[LoadQueue.scala 192:53:@38681.4]
  wire [1:0] _T_89764; // @[LoadQueue.scala 191:60:@38738.4]
  wire [1:0] _T_89765; // @[LoadQueue.scala 191:60:@38739.4]
  wire [2:0] _T_89766; // @[LoadQueue.scala 191:60:@38740.4]
  wire [2:0] _T_89767; // @[LoadQueue.scala 191:60:@38741.4]
  wire [2:0] _T_89768; // @[LoadQueue.scala 191:60:@38742.4]
  wire [2:0] _T_89769; // @[LoadQueue.scala 191:60:@38743.4]
  wire [3:0] _T_89770; // @[LoadQueue.scala 191:60:@38744.4]
  wire [3:0] _T_89771; // @[LoadQueue.scala 191:60:@38745.4]
  wire [3:0] _T_89772; // @[LoadQueue.scala 191:60:@38746.4]
  wire [3:0] _T_89773; // @[LoadQueue.scala 191:60:@38747.4]
  wire [3:0] _T_89774; // @[LoadQueue.scala 191:60:@38748.4]
  wire [3:0] _T_89775; // @[LoadQueue.scala 191:60:@38749.4]
  wire [3:0] _T_89776; // @[LoadQueue.scala 191:60:@38750.4]
  wire [3:0] _T_89777; // @[LoadQueue.scala 191:60:@38751.4]
  wire  _T_89780; // @[LoadQueue.scala 192:43:@38753.4]
  wire  _T_89781; // @[LoadQueue.scala 192:43:@38754.4]
  wire  _T_89782; // @[LoadQueue.scala 192:43:@38755.4]
  wire  _T_89783; // @[LoadQueue.scala 192:43:@38756.4]
  wire  _T_89784; // @[LoadQueue.scala 192:43:@38757.4]
  wire  _T_89785; // @[LoadQueue.scala 192:43:@38758.4]
  wire  _T_89786; // @[LoadQueue.scala 192:43:@38759.4]
  wire  _T_89787; // @[LoadQueue.scala 192:43:@38760.4]
  wire  _T_89788; // @[LoadQueue.scala 192:43:@38761.4]
  wire  _T_89789; // @[LoadQueue.scala 192:43:@38762.4]
  wire  _T_89790; // @[LoadQueue.scala 192:43:@38763.4]
  wire  _T_89791; // @[LoadQueue.scala 192:43:@38764.4]
  wire  _T_89792; // @[LoadQueue.scala 192:43:@38765.4]
  wire  _T_89793; // @[LoadQueue.scala 192:43:@38766.4]
  wire  _T_89794; // @[LoadQueue.scala 192:43:@38767.4]
  wire  _GEN_1590; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1591; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1592; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1593; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1594; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1595; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1596; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1597; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1598; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1599; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1600; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1601; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1602; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1603; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1604; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1605; // @[LoadQueue.scala 193:43:@38769.6]
  wire  _GEN_1607; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1608; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1609; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1610; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1611; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1612; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1613; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1614; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1615; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1616; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1617; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1618; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1619; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1620; // @[LoadQueue.scala 194:31:@38770.6]
  wire  _GEN_1621; // @[LoadQueue.scala 194:31:@38770.6]
  wire [31:0] _GEN_1623; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1624; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1625; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1626; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1627; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1628; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1629; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1630; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1631; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1632; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1633; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1634; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1635; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1636; // @[LoadQueue.scala 195:31:@38771.6]
  wire [31:0] _GEN_1637; // @[LoadQueue.scala 195:31:@38771.6]
  wire  lastConflict_11_0; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_1; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_2; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_3; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_4; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_5; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_6; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_7; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_8; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_9; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_10; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_11; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_12; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_13; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_14; // @[LoadQueue.scala 192:53:@38768.4]
  wire  lastConflict_11_15; // @[LoadQueue.scala 192:53:@38768.4]
  wire  canBypass_11; // @[LoadQueue.scala 192:53:@38768.4]
  wire [31:0] bypassVal_11; // @[LoadQueue.scala 192:53:@38768.4]
  wire [1:0] _T_89900; // @[LoadQueue.scala 191:60:@38825.4]
  wire [1:0] _T_89901; // @[LoadQueue.scala 191:60:@38826.4]
  wire [2:0] _T_89902; // @[LoadQueue.scala 191:60:@38827.4]
  wire [2:0] _T_89903; // @[LoadQueue.scala 191:60:@38828.4]
  wire [2:0] _T_89904; // @[LoadQueue.scala 191:60:@38829.4]
  wire [2:0] _T_89905; // @[LoadQueue.scala 191:60:@38830.4]
  wire [3:0] _T_89906; // @[LoadQueue.scala 191:60:@38831.4]
  wire [3:0] _T_89907; // @[LoadQueue.scala 191:60:@38832.4]
  wire [3:0] _T_89908; // @[LoadQueue.scala 191:60:@38833.4]
  wire [3:0] _T_89909; // @[LoadQueue.scala 191:60:@38834.4]
  wire [3:0] _T_89910; // @[LoadQueue.scala 191:60:@38835.4]
  wire [3:0] _T_89911; // @[LoadQueue.scala 191:60:@38836.4]
  wire [3:0] _T_89912; // @[LoadQueue.scala 191:60:@38837.4]
  wire [3:0] _T_89913; // @[LoadQueue.scala 191:60:@38838.4]
  wire  _T_89916; // @[LoadQueue.scala 192:43:@38840.4]
  wire  _T_89917; // @[LoadQueue.scala 192:43:@38841.4]
  wire  _T_89918; // @[LoadQueue.scala 192:43:@38842.4]
  wire  _T_89919; // @[LoadQueue.scala 192:43:@38843.4]
  wire  _T_89920; // @[LoadQueue.scala 192:43:@38844.4]
  wire  _T_89921; // @[LoadQueue.scala 192:43:@38845.4]
  wire  _T_89922; // @[LoadQueue.scala 192:43:@38846.4]
  wire  _T_89923; // @[LoadQueue.scala 192:43:@38847.4]
  wire  _T_89924; // @[LoadQueue.scala 192:43:@38848.4]
  wire  _T_89925; // @[LoadQueue.scala 192:43:@38849.4]
  wire  _T_89926; // @[LoadQueue.scala 192:43:@38850.4]
  wire  _T_89927; // @[LoadQueue.scala 192:43:@38851.4]
  wire  _T_89928; // @[LoadQueue.scala 192:43:@38852.4]
  wire  _T_89929; // @[LoadQueue.scala 192:43:@38853.4]
  wire  _T_89930; // @[LoadQueue.scala 192:43:@38854.4]
  wire  _GEN_1656; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1657; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1658; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1659; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1660; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1661; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1662; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1663; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1664; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1665; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1666; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1667; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1668; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1669; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1670; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1671; // @[LoadQueue.scala 193:43:@38856.6]
  wire  _GEN_1673; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1674; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1675; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1676; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1677; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1678; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1679; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1680; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1681; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1682; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1683; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1684; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1685; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1686; // @[LoadQueue.scala 194:31:@38857.6]
  wire  _GEN_1687; // @[LoadQueue.scala 194:31:@38857.6]
  wire [31:0] _GEN_1689; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1690; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1691; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1692; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1693; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1694; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1695; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1696; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1697; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1698; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1699; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1700; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1701; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1702; // @[LoadQueue.scala 195:31:@38858.6]
  wire [31:0] _GEN_1703; // @[LoadQueue.scala 195:31:@38858.6]
  wire  lastConflict_12_0; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_1; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_2; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_3; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_4; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_5; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_6; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_7; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_8; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_9; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_10; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_11; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_12; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_13; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_14; // @[LoadQueue.scala 192:53:@38855.4]
  wire  lastConflict_12_15; // @[LoadQueue.scala 192:53:@38855.4]
  wire  canBypass_12; // @[LoadQueue.scala 192:53:@38855.4]
  wire [31:0] bypassVal_12; // @[LoadQueue.scala 192:53:@38855.4]
  wire [1:0] _T_90036; // @[LoadQueue.scala 191:60:@38912.4]
  wire [1:0] _T_90037; // @[LoadQueue.scala 191:60:@38913.4]
  wire [2:0] _T_90038; // @[LoadQueue.scala 191:60:@38914.4]
  wire [2:0] _T_90039; // @[LoadQueue.scala 191:60:@38915.4]
  wire [2:0] _T_90040; // @[LoadQueue.scala 191:60:@38916.4]
  wire [2:0] _T_90041; // @[LoadQueue.scala 191:60:@38917.4]
  wire [3:0] _T_90042; // @[LoadQueue.scala 191:60:@38918.4]
  wire [3:0] _T_90043; // @[LoadQueue.scala 191:60:@38919.4]
  wire [3:0] _T_90044; // @[LoadQueue.scala 191:60:@38920.4]
  wire [3:0] _T_90045; // @[LoadQueue.scala 191:60:@38921.4]
  wire [3:0] _T_90046; // @[LoadQueue.scala 191:60:@38922.4]
  wire [3:0] _T_90047; // @[LoadQueue.scala 191:60:@38923.4]
  wire [3:0] _T_90048; // @[LoadQueue.scala 191:60:@38924.4]
  wire [3:0] _T_90049; // @[LoadQueue.scala 191:60:@38925.4]
  wire  _T_90052; // @[LoadQueue.scala 192:43:@38927.4]
  wire  _T_90053; // @[LoadQueue.scala 192:43:@38928.4]
  wire  _T_90054; // @[LoadQueue.scala 192:43:@38929.4]
  wire  _T_90055; // @[LoadQueue.scala 192:43:@38930.4]
  wire  _T_90056; // @[LoadQueue.scala 192:43:@38931.4]
  wire  _T_90057; // @[LoadQueue.scala 192:43:@38932.4]
  wire  _T_90058; // @[LoadQueue.scala 192:43:@38933.4]
  wire  _T_90059; // @[LoadQueue.scala 192:43:@38934.4]
  wire  _T_90060; // @[LoadQueue.scala 192:43:@38935.4]
  wire  _T_90061; // @[LoadQueue.scala 192:43:@38936.4]
  wire  _T_90062; // @[LoadQueue.scala 192:43:@38937.4]
  wire  _T_90063; // @[LoadQueue.scala 192:43:@38938.4]
  wire  _T_90064; // @[LoadQueue.scala 192:43:@38939.4]
  wire  _T_90065; // @[LoadQueue.scala 192:43:@38940.4]
  wire  _T_90066; // @[LoadQueue.scala 192:43:@38941.4]
  wire  _GEN_1722; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1723; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1724; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1725; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1726; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1727; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1728; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1729; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1730; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1731; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1732; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1733; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1734; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1735; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1736; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1737; // @[LoadQueue.scala 193:43:@38943.6]
  wire  _GEN_1739; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1740; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1741; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1742; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1743; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1744; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1745; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1746; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1747; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1748; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1749; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1750; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1751; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1752; // @[LoadQueue.scala 194:31:@38944.6]
  wire  _GEN_1753; // @[LoadQueue.scala 194:31:@38944.6]
  wire [31:0] _GEN_1755; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1756; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1757; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1758; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1759; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1760; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1761; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1762; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1763; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1764; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1765; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1766; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1767; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1768; // @[LoadQueue.scala 195:31:@38945.6]
  wire [31:0] _GEN_1769; // @[LoadQueue.scala 195:31:@38945.6]
  wire  lastConflict_13_0; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_1; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_2; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_3; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_4; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_5; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_6; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_7; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_8; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_9; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_10; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_11; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_12; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_13; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_14; // @[LoadQueue.scala 192:53:@38942.4]
  wire  lastConflict_13_15; // @[LoadQueue.scala 192:53:@38942.4]
  wire  canBypass_13; // @[LoadQueue.scala 192:53:@38942.4]
  wire [31:0] bypassVal_13; // @[LoadQueue.scala 192:53:@38942.4]
  wire [1:0] _T_90172; // @[LoadQueue.scala 191:60:@38999.4]
  wire [1:0] _T_90173; // @[LoadQueue.scala 191:60:@39000.4]
  wire [2:0] _T_90174; // @[LoadQueue.scala 191:60:@39001.4]
  wire [2:0] _T_90175; // @[LoadQueue.scala 191:60:@39002.4]
  wire [2:0] _T_90176; // @[LoadQueue.scala 191:60:@39003.4]
  wire [2:0] _T_90177; // @[LoadQueue.scala 191:60:@39004.4]
  wire [3:0] _T_90178; // @[LoadQueue.scala 191:60:@39005.4]
  wire [3:0] _T_90179; // @[LoadQueue.scala 191:60:@39006.4]
  wire [3:0] _T_90180; // @[LoadQueue.scala 191:60:@39007.4]
  wire [3:0] _T_90181; // @[LoadQueue.scala 191:60:@39008.4]
  wire [3:0] _T_90182; // @[LoadQueue.scala 191:60:@39009.4]
  wire [3:0] _T_90183; // @[LoadQueue.scala 191:60:@39010.4]
  wire [3:0] _T_90184; // @[LoadQueue.scala 191:60:@39011.4]
  wire [3:0] _T_90185; // @[LoadQueue.scala 191:60:@39012.4]
  wire  _T_90188; // @[LoadQueue.scala 192:43:@39014.4]
  wire  _T_90189; // @[LoadQueue.scala 192:43:@39015.4]
  wire  _T_90190; // @[LoadQueue.scala 192:43:@39016.4]
  wire  _T_90191; // @[LoadQueue.scala 192:43:@39017.4]
  wire  _T_90192; // @[LoadQueue.scala 192:43:@39018.4]
  wire  _T_90193; // @[LoadQueue.scala 192:43:@39019.4]
  wire  _T_90194; // @[LoadQueue.scala 192:43:@39020.4]
  wire  _T_90195; // @[LoadQueue.scala 192:43:@39021.4]
  wire  _T_90196; // @[LoadQueue.scala 192:43:@39022.4]
  wire  _T_90197; // @[LoadQueue.scala 192:43:@39023.4]
  wire  _T_90198; // @[LoadQueue.scala 192:43:@39024.4]
  wire  _T_90199; // @[LoadQueue.scala 192:43:@39025.4]
  wire  _T_90200; // @[LoadQueue.scala 192:43:@39026.4]
  wire  _T_90201; // @[LoadQueue.scala 192:43:@39027.4]
  wire  _T_90202; // @[LoadQueue.scala 192:43:@39028.4]
  wire  _GEN_1788; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1789; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1790; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1791; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1792; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1793; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1794; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1795; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1796; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1797; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1798; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1799; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1800; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1801; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1802; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1803; // @[LoadQueue.scala 193:43:@39030.6]
  wire  _GEN_1805; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1806; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1807; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1808; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1809; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1810; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1811; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1812; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1813; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1814; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1815; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1816; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1817; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1818; // @[LoadQueue.scala 194:31:@39031.6]
  wire  _GEN_1819; // @[LoadQueue.scala 194:31:@39031.6]
  wire [31:0] _GEN_1821; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1822; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1823; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1824; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1825; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1826; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1827; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1828; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1829; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1830; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1831; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1832; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1833; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1834; // @[LoadQueue.scala 195:31:@39032.6]
  wire [31:0] _GEN_1835; // @[LoadQueue.scala 195:31:@39032.6]
  wire  lastConflict_14_0; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_1; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_2; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_3; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_4; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_5; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_6; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_7; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_8; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_9; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_10; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_11; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_12; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_13; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_14; // @[LoadQueue.scala 192:53:@39029.4]
  wire  lastConflict_14_15; // @[LoadQueue.scala 192:53:@39029.4]
  wire  canBypass_14; // @[LoadQueue.scala 192:53:@39029.4]
  wire [31:0] bypassVal_14; // @[LoadQueue.scala 192:53:@39029.4]
  wire [1:0] _T_90308; // @[LoadQueue.scala 191:60:@39086.4]
  wire [1:0] _T_90309; // @[LoadQueue.scala 191:60:@39087.4]
  wire [2:0] _T_90310; // @[LoadQueue.scala 191:60:@39088.4]
  wire [2:0] _T_90311; // @[LoadQueue.scala 191:60:@39089.4]
  wire [2:0] _T_90312; // @[LoadQueue.scala 191:60:@39090.4]
  wire [2:0] _T_90313; // @[LoadQueue.scala 191:60:@39091.4]
  wire [3:0] _T_90314; // @[LoadQueue.scala 191:60:@39092.4]
  wire [3:0] _T_90315; // @[LoadQueue.scala 191:60:@39093.4]
  wire [3:0] _T_90316; // @[LoadQueue.scala 191:60:@39094.4]
  wire [3:0] _T_90317; // @[LoadQueue.scala 191:60:@39095.4]
  wire [3:0] _T_90318; // @[LoadQueue.scala 191:60:@39096.4]
  wire [3:0] _T_90319; // @[LoadQueue.scala 191:60:@39097.4]
  wire [3:0] _T_90320; // @[LoadQueue.scala 191:60:@39098.4]
  wire [3:0] _T_90321; // @[LoadQueue.scala 191:60:@39099.4]
  wire  _T_90324; // @[LoadQueue.scala 192:43:@39101.4]
  wire  _T_90325; // @[LoadQueue.scala 192:43:@39102.4]
  wire  _T_90326; // @[LoadQueue.scala 192:43:@39103.4]
  wire  _T_90327; // @[LoadQueue.scala 192:43:@39104.4]
  wire  _T_90328; // @[LoadQueue.scala 192:43:@39105.4]
  wire  _T_90329; // @[LoadQueue.scala 192:43:@39106.4]
  wire  _T_90330; // @[LoadQueue.scala 192:43:@39107.4]
  wire  _T_90331; // @[LoadQueue.scala 192:43:@39108.4]
  wire  _T_90332; // @[LoadQueue.scala 192:43:@39109.4]
  wire  _T_90333; // @[LoadQueue.scala 192:43:@39110.4]
  wire  _T_90334; // @[LoadQueue.scala 192:43:@39111.4]
  wire  _T_90335; // @[LoadQueue.scala 192:43:@39112.4]
  wire  _T_90336; // @[LoadQueue.scala 192:43:@39113.4]
  wire  _T_90337; // @[LoadQueue.scala 192:43:@39114.4]
  wire  _T_90338; // @[LoadQueue.scala 192:43:@39115.4]
  wire  _GEN_1854; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1855; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1856; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1857; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1858; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1859; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1860; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1861; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1862; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1863; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1864; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1865; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1866; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1867; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1868; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1869; // @[LoadQueue.scala 193:43:@39117.6]
  wire  _GEN_1871; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1872; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1873; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1874; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1875; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1876; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1877; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1878; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1879; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1880; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1881; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1882; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1883; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1884; // @[LoadQueue.scala 194:31:@39118.6]
  wire  _GEN_1885; // @[LoadQueue.scala 194:31:@39118.6]
  wire [31:0] _GEN_1887; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1888; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1889; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1890; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1891; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1892; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1893; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1894; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1895; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1896; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1897; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1898; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1899; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1900; // @[LoadQueue.scala 195:31:@39119.6]
  wire [31:0] _GEN_1901; // @[LoadQueue.scala 195:31:@39119.6]
  wire  lastConflict_15_0; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_1; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_2; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_3; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_4; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_5; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_6; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_7; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_8; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_9; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_10; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_11; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_12; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_13; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_14; // @[LoadQueue.scala 192:53:@39116.4]
  wire  lastConflict_15_15; // @[LoadQueue.scala 192:53:@39116.4]
  wire  canBypass_15; // @[LoadQueue.scala 192:53:@39116.4]
  wire [31:0] bypassVal_15; // @[LoadQueue.scala 192:53:@39116.4]
  wire [15:0] _T_90398; // @[OneHot.scala 52:12:@39124.4]
  wire  _T_90400; // @[util.scala 33:60:@39126.4]
  wire  _T_90401; // @[util.scala 33:60:@39127.4]
  wire  _T_90402; // @[util.scala 33:60:@39128.4]
  wire  _T_90403; // @[util.scala 33:60:@39129.4]
  wire  _T_90404; // @[util.scala 33:60:@39130.4]
  wire  _T_90405; // @[util.scala 33:60:@39131.4]
  wire  _T_90406; // @[util.scala 33:60:@39132.4]
  wire  _T_90407; // @[util.scala 33:60:@39133.4]
  wire  _T_90408; // @[util.scala 33:60:@39134.4]
  wire  _T_90409; // @[util.scala 33:60:@39135.4]
  wire  _T_90410; // @[util.scala 33:60:@39136.4]
  wire  _T_90411; // @[util.scala 33:60:@39137.4]
  wire  _T_90412; // @[util.scala 33:60:@39138.4]
  wire  _T_90413; // @[util.scala 33:60:@39139.4]
  wire  _T_90414; // @[util.scala 33:60:@39140.4]
  wire  _T_90415; // @[util.scala 33:60:@39141.4]
  wire  _T_93512; // @[LoadQueue.scala 229:41:@41664.4]
  wire  _T_93513; // @[LoadQueue.scala 229:38:@41665.4]
  wire  _T_93515; // @[LoadQueue.scala 230:12:@41667.6]
  reg  prevPriorityRequest_15; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_739;
  wire  _T_93517; // @[LoadQueue.scala 230:46:@41668.6]
  wire  _T_93518; // @[LoadQueue.scala 230:43:@41669.6]
  wire  _T_93520; // @[LoadQueue.scala 230:84:@41670.6]
  wire  _T_93521; // @[LoadQueue.scala 230:81:@41671.6]
  wire  _T_93524; // @[LoadQueue.scala 233:86:@41674.8]
  wire  _T_93525; // @[LoadQueue.scala 233:86:@41675.8]
  wire  _T_93526; // @[LoadQueue.scala 233:86:@41676.8]
  wire  _T_93527; // @[LoadQueue.scala 233:86:@41677.8]
  wire  _T_93528; // @[LoadQueue.scala 233:86:@41678.8]
  wire  _T_93529; // @[LoadQueue.scala 233:86:@41679.8]
  wire  _T_93530; // @[LoadQueue.scala 233:86:@41680.8]
  wire  _T_93531; // @[LoadQueue.scala 233:86:@41681.8]
  wire  _T_93532; // @[LoadQueue.scala 233:86:@41682.8]
  wire  _T_93533; // @[LoadQueue.scala 233:86:@41683.8]
  wire  _T_93534; // @[LoadQueue.scala 233:86:@41684.8]
  wire  _T_93535; // @[LoadQueue.scala 233:86:@41685.8]
  wire  _T_93536; // @[LoadQueue.scala 233:86:@41686.8]
  wire  _T_93537; // @[LoadQueue.scala 233:86:@41687.8]
  wire  _T_93538; // @[LoadQueue.scala 233:86:@41688.8]
  wire  _T_93540; // @[LoadQueue.scala 233:38:@41689.8]
  wire  _T_93559; // @[LoadQueue.scala 234:11:@41706.8]
  wire  _T_93560; // @[LoadQueue.scala 233:103:@41707.8]
  wire  _GEN_2028; // @[LoadQueue.scala 230:110:@41672.6]
  wire  loadRequest_15; // @[LoadQueue.scala 229:71:@41666.4]
  wire [15:0] _T_90456; // @[Mux.scala 31:69:@39159.4]
  wire  _T_93428; // @[LoadQueue.scala 229:41:@41582.4]
  wire  _T_93429; // @[LoadQueue.scala 229:38:@41583.4]
  wire  _T_93431; // @[LoadQueue.scala 230:12:@41585.6]
  reg  prevPriorityRequest_14; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_740;
  wire  _T_93433; // @[LoadQueue.scala 230:46:@41586.6]
  wire  _T_93434; // @[LoadQueue.scala 230:43:@41587.6]
  wire  _T_93436; // @[LoadQueue.scala 230:84:@41588.6]
  wire  _T_93437; // @[LoadQueue.scala 230:81:@41589.6]
  wire  _T_93440; // @[LoadQueue.scala 233:86:@41592.8]
  wire  _T_93441; // @[LoadQueue.scala 233:86:@41593.8]
  wire  _T_93442; // @[LoadQueue.scala 233:86:@41594.8]
  wire  _T_93443; // @[LoadQueue.scala 233:86:@41595.8]
  wire  _T_93444; // @[LoadQueue.scala 233:86:@41596.8]
  wire  _T_93445; // @[LoadQueue.scala 233:86:@41597.8]
  wire  _T_93446; // @[LoadQueue.scala 233:86:@41598.8]
  wire  _T_93447; // @[LoadQueue.scala 233:86:@41599.8]
  wire  _T_93448; // @[LoadQueue.scala 233:86:@41600.8]
  wire  _T_93449; // @[LoadQueue.scala 233:86:@41601.8]
  wire  _T_93450; // @[LoadQueue.scala 233:86:@41602.8]
  wire  _T_93451; // @[LoadQueue.scala 233:86:@41603.8]
  wire  _T_93452; // @[LoadQueue.scala 233:86:@41604.8]
  wire  _T_93453; // @[LoadQueue.scala 233:86:@41605.8]
  wire  _T_93454; // @[LoadQueue.scala 233:86:@41606.8]
  wire  _T_93456; // @[LoadQueue.scala 233:38:@41607.8]
  wire  _T_93475; // @[LoadQueue.scala 234:11:@41624.8]
  wire  _T_93476; // @[LoadQueue.scala 233:103:@41625.8]
  wire  _GEN_2024; // @[LoadQueue.scala 230:110:@41590.6]
  wire  loadRequest_14; // @[LoadQueue.scala 229:71:@41584.4]
  wire [15:0] _T_90457; // @[Mux.scala 31:69:@39160.4]
  wire  _T_93344; // @[LoadQueue.scala 229:41:@41500.4]
  wire  _T_93345; // @[LoadQueue.scala 229:38:@41501.4]
  wire  _T_93347; // @[LoadQueue.scala 230:12:@41503.6]
  reg  prevPriorityRequest_13; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_741;
  wire  _T_93349; // @[LoadQueue.scala 230:46:@41504.6]
  wire  _T_93350; // @[LoadQueue.scala 230:43:@41505.6]
  wire  _T_93352; // @[LoadQueue.scala 230:84:@41506.6]
  wire  _T_93353; // @[LoadQueue.scala 230:81:@41507.6]
  wire  _T_93356; // @[LoadQueue.scala 233:86:@41510.8]
  wire  _T_93357; // @[LoadQueue.scala 233:86:@41511.8]
  wire  _T_93358; // @[LoadQueue.scala 233:86:@41512.8]
  wire  _T_93359; // @[LoadQueue.scala 233:86:@41513.8]
  wire  _T_93360; // @[LoadQueue.scala 233:86:@41514.8]
  wire  _T_93361; // @[LoadQueue.scala 233:86:@41515.8]
  wire  _T_93362; // @[LoadQueue.scala 233:86:@41516.8]
  wire  _T_93363; // @[LoadQueue.scala 233:86:@41517.8]
  wire  _T_93364; // @[LoadQueue.scala 233:86:@41518.8]
  wire  _T_93365; // @[LoadQueue.scala 233:86:@41519.8]
  wire  _T_93366; // @[LoadQueue.scala 233:86:@41520.8]
  wire  _T_93367; // @[LoadQueue.scala 233:86:@41521.8]
  wire  _T_93368; // @[LoadQueue.scala 233:86:@41522.8]
  wire  _T_93369; // @[LoadQueue.scala 233:86:@41523.8]
  wire  _T_93370; // @[LoadQueue.scala 233:86:@41524.8]
  wire  _T_93372; // @[LoadQueue.scala 233:38:@41525.8]
  wire  _T_93391; // @[LoadQueue.scala 234:11:@41542.8]
  wire  _T_93392; // @[LoadQueue.scala 233:103:@41543.8]
  wire  _GEN_2020; // @[LoadQueue.scala 230:110:@41508.6]
  wire  loadRequest_13; // @[LoadQueue.scala 229:71:@41502.4]
  wire [15:0] _T_90458; // @[Mux.scala 31:69:@39161.4]
  wire  _T_93260; // @[LoadQueue.scala 229:41:@41418.4]
  wire  _T_93261; // @[LoadQueue.scala 229:38:@41419.4]
  wire  _T_93263; // @[LoadQueue.scala 230:12:@41421.6]
  reg  prevPriorityRequest_12; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_742;
  wire  _T_93265; // @[LoadQueue.scala 230:46:@41422.6]
  wire  _T_93266; // @[LoadQueue.scala 230:43:@41423.6]
  wire  _T_93268; // @[LoadQueue.scala 230:84:@41424.6]
  wire  _T_93269; // @[LoadQueue.scala 230:81:@41425.6]
  wire  _T_93272; // @[LoadQueue.scala 233:86:@41428.8]
  wire  _T_93273; // @[LoadQueue.scala 233:86:@41429.8]
  wire  _T_93274; // @[LoadQueue.scala 233:86:@41430.8]
  wire  _T_93275; // @[LoadQueue.scala 233:86:@41431.8]
  wire  _T_93276; // @[LoadQueue.scala 233:86:@41432.8]
  wire  _T_93277; // @[LoadQueue.scala 233:86:@41433.8]
  wire  _T_93278; // @[LoadQueue.scala 233:86:@41434.8]
  wire  _T_93279; // @[LoadQueue.scala 233:86:@41435.8]
  wire  _T_93280; // @[LoadQueue.scala 233:86:@41436.8]
  wire  _T_93281; // @[LoadQueue.scala 233:86:@41437.8]
  wire  _T_93282; // @[LoadQueue.scala 233:86:@41438.8]
  wire  _T_93283; // @[LoadQueue.scala 233:86:@41439.8]
  wire  _T_93284; // @[LoadQueue.scala 233:86:@41440.8]
  wire  _T_93285; // @[LoadQueue.scala 233:86:@41441.8]
  wire  _T_93286; // @[LoadQueue.scala 233:86:@41442.8]
  wire  _T_93288; // @[LoadQueue.scala 233:38:@41443.8]
  wire  _T_93307; // @[LoadQueue.scala 234:11:@41460.8]
  wire  _T_93308; // @[LoadQueue.scala 233:103:@41461.8]
  wire  _GEN_2016; // @[LoadQueue.scala 230:110:@41426.6]
  wire  loadRequest_12; // @[LoadQueue.scala 229:71:@41420.4]
  wire [15:0] _T_90459; // @[Mux.scala 31:69:@39162.4]
  wire  _T_93176; // @[LoadQueue.scala 229:41:@41336.4]
  wire  _T_93177; // @[LoadQueue.scala 229:38:@41337.4]
  wire  _T_93179; // @[LoadQueue.scala 230:12:@41339.6]
  reg  prevPriorityRequest_11; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_743;
  wire  _T_93181; // @[LoadQueue.scala 230:46:@41340.6]
  wire  _T_93182; // @[LoadQueue.scala 230:43:@41341.6]
  wire  _T_93184; // @[LoadQueue.scala 230:84:@41342.6]
  wire  _T_93185; // @[LoadQueue.scala 230:81:@41343.6]
  wire  _T_93188; // @[LoadQueue.scala 233:86:@41346.8]
  wire  _T_93189; // @[LoadQueue.scala 233:86:@41347.8]
  wire  _T_93190; // @[LoadQueue.scala 233:86:@41348.8]
  wire  _T_93191; // @[LoadQueue.scala 233:86:@41349.8]
  wire  _T_93192; // @[LoadQueue.scala 233:86:@41350.8]
  wire  _T_93193; // @[LoadQueue.scala 233:86:@41351.8]
  wire  _T_93194; // @[LoadQueue.scala 233:86:@41352.8]
  wire  _T_93195; // @[LoadQueue.scala 233:86:@41353.8]
  wire  _T_93196; // @[LoadQueue.scala 233:86:@41354.8]
  wire  _T_93197; // @[LoadQueue.scala 233:86:@41355.8]
  wire  _T_93198; // @[LoadQueue.scala 233:86:@41356.8]
  wire  _T_93199; // @[LoadQueue.scala 233:86:@41357.8]
  wire  _T_93200; // @[LoadQueue.scala 233:86:@41358.8]
  wire  _T_93201; // @[LoadQueue.scala 233:86:@41359.8]
  wire  _T_93202; // @[LoadQueue.scala 233:86:@41360.8]
  wire  _T_93204; // @[LoadQueue.scala 233:38:@41361.8]
  wire  _T_93223; // @[LoadQueue.scala 234:11:@41378.8]
  wire  _T_93224; // @[LoadQueue.scala 233:103:@41379.8]
  wire  _GEN_2012; // @[LoadQueue.scala 230:110:@41344.6]
  wire  loadRequest_11; // @[LoadQueue.scala 229:71:@41338.4]
  wire [15:0] _T_90460; // @[Mux.scala 31:69:@39163.4]
  wire  _T_93092; // @[LoadQueue.scala 229:41:@41254.4]
  wire  _T_93093; // @[LoadQueue.scala 229:38:@41255.4]
  wire  _T_93095; // @[LoadQueue.scala 230:12:@41257.6]
  reg  prevPriorityRequest_10; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_744;
  wire  _T_93097; // @[LoadQueue.scala 230:46:@41258.6]
  wire  _T_93098; // @[LoadQueue.scala 230:43:@41259.6]
  wire  _T_93100; // @[LoadQueue.scala 230:84:@41260.6]
  wire  _T_93101; // @[LoadQueue.scala 230:81:@41261.6]
  wire  _T_93104; // @[LoadQueue.scala 233:86:@41264.8]
  wire  _T_93105; // @[LoadQueue.scala 233:86:@41265.8]
  wire  _T_93106; // @[LoadQueue.scala 233:86:@41266.8]
  wire  _T_93107; // @[LoadQueue.scala 233:86:@41267.8]
  wire  _T_93108; // @[LoadQueue.scala 233:86:@41268.8]
  wire  _T_93109; // @[LoadQueue.scala 233:86:@41269.8]
  wire  _T_93110; // @[LoadQueue.scala 233:86:@41270.8]
  wire  _T_93111; // @[LoadQueue.scala 233:86:@41271.8]
  wire  _T_93112; // @[LoadQueue.scala 233:86:@41272.8]
  wire  _T_93113; // @[LoadQueue.scala 233:86:@41273.8]
  wire  _T_93114; // @[LoadQueue.scala 233:86:@41274.8]
  wire  _T_93115; // @[LoadQueue.scala 233:86:@41275.8]
  wire  _T_93116; // @[LoadQueue.scala 233:86:@41276.8]
  wire  _T_93117; // @[LoadQueue.scala 233:86:@41277.8]
  wire  _T_93118; // @[LoadQueue.scala 233:86:@41278.8]
  wire  _T_93120; // @[LoadQueue.scala 233:38:@41279.8]
  wire  _T_93139; // @[LoadQueue.scala 234:11:@41296.8]
  wire  _T_93140; // @[LoadQueue.scala 233:103:@41297.8]
  wire  _GEN_2008; // @[LoadQueue.scala 230:110:@41262.6]
  wire  loadRequest_10; // @[LoadQueue.scala 229:71:@41256.4]
  wire [15:0] _T_90461; // @[Mux.scala 31:69:@39164.4]
  wire  _T_93008; // @[LoadQueue.scala 229:41:@41172.4]
  wire  _T_93009; // @[LoadQueue.scala 229:38:@41173.4]
  wire  _T_93011; // @[LoadQueue.scala 230:12:@41175.6]
  reg  prevPriorityRequest_9; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_745;
  wire  _T_93013; // @[LoadQueue.scala 230:46:@41176.6]
  wire  _T_93014; // @[LoadQueue.scala 230:43:@41177.6]
  wire  _T_93016; // @[LoadQueue.scala 230:84:@41178.6]
  wire  _T_93017; // @[LoadQueue.scala 230:81:@41179.6]
  wire  _T_93020; // @[LoadQueue.scala 233:86:@41182.8]
  wire  _T_93021; // @[LoadQueue.scala 233:86:@41183.8]
  wire  _T_93022; // @[LoadQueue.scala 233:86:@41184.8]
  wire  _T_93023; // @[LoadQueue.scala 233:86:@41185.8]
  wire  _T_93024; // @[LoadQueue.scala 233:86:@41186.8]
  wire  _T_93025; // @[LoadQueue.scala 233:86:@41187.8]
  wire  _T_93026; // @[LoadQueue.scala 233:86:@41188.8]
  wire  _T_93027; // @[LoadQueue.scala 233:86:@41189.8]
  wire  _T_93028; // @[LoadQueue.scala 233:86:@41190.8]
  wire  _T_93029; // @[LoadQueue.scala 233:86:@41191.8]
  wire  _T_93030; // @[LoadQueue.scala 233:86:@41192.8]
  wire  _T_93031; // @[LoadQueue.scala 233:86:@41193.8]
  wire  _T_93032; // @[LoadQueue.scala 233:86:@41194.8]
  wire  _T_93033; // @[LoadQueue.scala 233:86:@41195.8]
  wire  _T_93034; // @[LoadQueue.scala 233:86:@41196.8]
  wire  _T_93036; // @[LoadQueue.scala 233:38:@41197.8]
  wire  _T_93055; // @[LoadQueue.scala 234:11:@41214.8]
  wire  _T_93056; // @[LoadQueue.scala 233:103:@41215.8]
  wire  _GEN_2004; // @[LoadQueue.scala 230:110:@41180.6]
  wire  loadRequest_9; // @[LoadQueue.scala 229:71:@41174.4]
  wire [15:0] _T_90462; // @[Mux.scala 31:69:@39165.4]
  wire  _T_92924; // @[LoadQueue.scala 229:41:@41090.4]
  wire  _T_92925; // @[LoadQueue.scala 229:38:@41091.4]
  wire  _T_92927; // @[LoadQueue.scala 230:12:@41093.6]
  reg  prevPriorityRequest_8; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_746;
  wire  _T_92929; // @[LoadQueue.scala 230:46:@41094.6]
  wire  _T_92930; // @[LoadQueue.scala 230:43:@41095.6]
  wire  _T_92932; // @[LoadQueue.scala 230:84:@41096.6]
  wire  _T_92933; // @[LoadQueue.scala 230:81:@41097.6]
  wire  _T_92936; // @[LoadQueue.scala 233:86:@41100.8]
  wire  _T_92937; // @[LoadQueue.scala 233:86:@41101.8]
  wire  _T_92938; // @[LoadQueue.scala 233:86:@41102.8]
  wire  _T_92939; // @[LoadQueue.scala 233:86:@41103.8]
  wire  _T_92940; // @[LoadQueue.scala 233:86:@41104.8]
  wire  _T_92941; // @[LoadQueue.scala 233:86:@41105.8]
  wire  _T_92942; // @[LoadQueue.scala 233:86:@41106.8]
  wire  _T_92943; // @[LoadQueue.scala 233:86:@41107.8]
  wire  _T_92944; // @[LoadQueue.scala 233:86:@41108.8]
  wire  _T_92945; // @[LoadQueue.scala 233:86:@41109.8]
  wire  _T_92946; // @[LoadQueue.scala 233:86:@41110.8]
  wire  _T_92947; // @[LoadQueue.scala 233:86:@41111.8]
  wire  _T_92948; // @[LoadQueue.scala 233:86:@41112.8]
  wire  _T_92949; // @[LoadQueue.scala 233:86:@41113.8]
  wire  _T_92950; // @[LoadQueue.scala 233:86:@41114.8]
  wire  _T_92952; // @[LoadQueue.scala 233:38:@41115.8]
  wire  _T_92971; // @[LoadQueue.scala 234:11:@41132.8]
  wire  _T_92972; // @[LoadQueue.scala 233:103:@41133.8]
  wire  _GEN_2000; // @[LoadQueue.scala 230:110:@41098.6]
  wire  loadRequest_8; // @[LoadQueue.scala 229:71:@41092.4]
  wire [15:0] _T_90463; // @[Mux.scala 31:69:@39166.4]
  wire  _T_92840; // @[LoadQueue.scala 229:41:@41008.4]
  wire  _T_92841; // @[LoadQueue.scala 229:38:@41009.4]
  wire  _T_92843; // @[LoadQueue.scala 230:12:@41011.6]
  reg  prevPriorityRequest_7; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_747;
  wire  _T_92845; // @[LoadQueue.scala 230:46:@41012.6]
  wire  _T_92846; // @[LoadQueue.scala 230:43:@41013.6]
  wire  _T_92848; // @[LoadQueue.scala 230:84:@41014.6]
  wire  _T_92849; // @[LoadQueue.scala 230:81:@41015.6]
  wire  _T_92852; // @[LoadQueue.scala 233:86:@41018.8]
  wire  _T_92853; // @[LoadQueue.scala 233:86:@41019.8]
  wire  _T_92854; // @[LoadQueue.scala 233:86:@41020.8]
  wire  _T_92855; // @[LoadQueue.scala 233:86:@41021.8]
  wire  _T_92856; // @[LoadQueue.scala 233:86:@41022.8]
  wire  _T_92857; // @[LoadQueue.scala 233:86:@41023.8]
  wire  _T_92858; // @[LoadQueue.scala 233:86:@41024.8]
  wire  _T_92859; // @[LoadQueue.scala 233:86:@41025.8]
  wire  _T_92860; // @[LoadQueue.scala 233:86:@41026.8]
  wire  _T_92861; // @[LoadQueue.scala 233:86:@41027.8]
  wire  _T_92862; // @[LoadQueue.scala 233:86:@41028.8]
  wire  _T_92863; // @[LoadQueue.scala 233:86:@41029.8]
  wire  _T_92864; // @[LoadQueue.scala 233:86:@41030.8]
  wire  _T_92865; // @[LoadQueue.scala 233:86:@41031.8]
  wire  _T_92866; // @[LoadQueue.scala 233:86:@41032.8]
  wire  _T_92868; // @[LoadQueue.scala 233:38:@41033.8]
  wire  _T_92887; // @[LoadQueue.scala 234:11:@41050.8]
  wire  _T_92888; // @[LoadQueue.scala 233:103:@41051.8]
  wire  _GEN_1996; // @[LoadQueue.scala 230:110:@41016.6]
  wire  loadRequest_7; // @[LoadQueue.scala 229:71:@41010.4]
  wire [15:0] _T_90464; // @[Mux.scala 31:69:@39167.4]
  wire  _T_92756; // @[LoadQueue.scala 229:41:@40926.4]
  wire  _T_92757; // @[LoadQueue.scala 229:38:@40927.4]
  wire  _T_92759; // @[LoadQueue.scala 230:12:@40929.6]
  reg  prevPriorityRequest_6; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_748;
  wire  _T_92761; // @[LoadQueue.scala 230:46:@40930.6]
  wire  _T_92762; // @[LoadQueue.scala 230:43:@40931.6]
  wire  _T_92764; // @[LoadQueue.scala 230:84:@40932.6]
  wire  _T_92765; // @[LoadQueue.scala 230:81:@40933.6]
  wire  _T_92768; // @[LoadQueue.scala 233:86:@40936.8]
  wire  _T_92769; // @[LoadQueue.scala 233:86:@40937.8]
  wire  _T_92770; // @[LoadQueue.scala 233:86:@40938.8]
  wire  _T_92771; // @[LoadQueue.scala 233:86:@40939.8]
  wire  _T_92772; // @[LoadQueue.scala 233:86:@40940.8]
  wire  _T_92773; // @[LoadQueue.scala 233:86:@40941.8]
  wire  _T_92774; // @[LoadQueue.scala 233:86:@40942.8]
  wire  _T_92775; // @[LoadQueue.scala 233:86:@40943.8]
  wire  _T_92776; // @[LoadQueue.scala 233:86:@40944.8]
  wire  _T_92777; // @[LoadQueue.scala 233:86:@40945.8]
  wire  _T_92778; // @[LoadQueue.scala 233:86:@40946.8]
  wire  _T_92779; // @[LoadQueue.scala 233:86:@40947.8]
  wire  _T_92780; // @[LoadQueue.scala 233:86:@40948.8]
  wire  _T_92781; // @[LoadQueue.scala 233:86:@40949.8]
  wire  _T_92782; // @[LoadQueue.scala 233:86:@40950.8]
  wire  _T_92784; // @[LoadQueue.scala 233:38:@40951.8]
  wire  _T_92803; // @[LoadQueue.scala 234:11:@40968.8]
  wire  _T_92804; // @[LoadQueue.scala 233:103:@40969.8]
  wire  _GEN_1992; // @[LoadQueue.scala 230:110:@40934.6]
  wire  loadRequest_6; // @[LoadQueue.scala 229:71:@40928.4]
  wire [15:0] _T_90465; // @[Mux.scala 31:69:@39168.4]
  wire  _T_92672; // @[LoadQueue.scala 229:41:@40844.4]
  wire  _T_92673; // @[LoadQueue.scala 229:38:@40845.4]
  wire  _T_92675; // @[LoadQueue.scala 230:12:@40847.6]
  reg  prevPriorityRequest_5; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_749;
  wire  _T_92677; // @[LoadQueue.scala 230:46:@40848.6]
  wire  _T_92678; // @[LoadQueue.scala 230:43:@40849.6]
  wire  _T_92680; // @[LoadQueue.scala 230:84:@40850.6]
  wire  _T_92681; // @[LoadQueue.scala 230:81:@40851.6]
  wire  _T_92684; // @[LoadQueue.scala 233:86:@40854.8]
  wire  _T_92685; // @[LoadQueue.scala 233:86:@40855.8]
  wire  _T_92686; // @[LoadQueue.scala 233:86:@40856.8]
  wire  _T_92687; // @[LoadQueue.scala 233:86:@40857.8]
  wire  _T_92688; // @[LoadQueue.scala 233:86:@40858.8]
  wire  _T_92689; // @[LoadQueue.scala 233:86:@40859.8]
  wire  _T_92690; // @[LoadQueue.scala 233:86:@40860.8]
  wire  _T_92691; // @[LoadQueue.scala 233:86:@40861.8]
  wire  _T_92692; // @[LoadQueue.scala 233:86:@40862.8]
  wire  _T_92693; // @[LoadQueue.scala 233:86:@40863.8]
  wire  _T_92694; // @[LoadQueue.scala 233:86:@40864.8]
  wire  _T_92695; // @[LoadQueue.scala 233:86:@40865.8]
  wire  _T_92696; // @[LoadQueue.scala 233:86:@40866.8]
  wire  _T_92697; // @[LoadQueue.scala 233:86:@40867.8]
  wire  _T_92698; // @[LoadQueue.scala 233:86:@40868.8]
  wire  _T_92700; // @[LoadQueue.scala 233:38:@40869.8]
  wire  _T_92719; // @[LoadQueue.scala 234:11:@40886.8]
  wire  _T_92720; // @[LoadQueue.scala 233:103:@40887.8]
  wire  _GEN_1988; // @[LoadQueue.scala 230:110:@40852.6]
  wire  loadRequest_5; // @[LoadQueue.scala 229:71:@40846.4]
  wire [15:0] _T_90466; // @[Mux.scala 31:69:@39169.4]
  wire  _T_92588; // @[LoadQueue.scala 229:41:@40762.4]
  wire  _T_92589; // @[LoadQueue.scala 229:38:@40763.4]
  wire  _T_92591; // @[LoadQueue.scala 230:12:@40765.6]
  reg  prevPriorityRequest_4; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_750;
  wire  _T_92593; // @[LoadQueue.scala 230:46:@40766.6]
  wire  _T_92594; // @[LoadQueue.scala 230:43:@40767.6]
  wire  _T_92596; // @[LoadQueue.scala 230:84:@40768.6]
  wire  _T_92597; // @[LoadQueue.scala 230:81:@40769.6]
  wire  _T_92600; // @[LoadQueue.scala 233:86:@40772.8]
  wire  _T_92601; // @[LoadQueue.scala 233:86:@40773.8]
  wire  _T_92602; // @[LoadQueue.scala 233:86:@40774.8]
  wire  _T_92603; // @[LoadQueue.scala 233:86:@40775.8]
  wire  _T_92604; // @[LoadQueue.scala 233:86:@40776.8]
  wire  _T_92605; // @[LoadQueue.scala 233:86:@40777.8]
  wire  _T_92606; // @[LoadQueue.scala 233:86:@40778.8]
  wire  _T_92607; // @[LoadQueue.scala 233:86:@40779.8]
  wire  _T_92608; // @[LoadQueue.scala 233:86:@40780.8]
  wire  _T_92609; // @[LoadQueue.scala 233:86:@40781.8]
  wire  _T_92610; // @[LoadQueue.scala 233:86:@40782.8]
  wire  _T_92611; // @[LoadQueue.scala 233:86:@40783.8]
  wire  _T_92612; // @[LoadQueue.scala 233:86:@40784.8]
  wire  _T_92613; // @[LoadQueue.scala 233:86:@40785.8]
  wire  _T_92614; // @[LoadQueue.scala 233:86:@40786.8]
  wire  _T_92616; // @[LoadQueue.scala 233:38:@40787.8]
  wire  _T_92635; // @[LoadQueue.scala 234:11:@40804.8]
  wire  _T_92636; // @[LoadQueue.scala 233:103:@40805.8]
  wire  _GEN_1984; // @[LoadQueue.scala 230:110:@40770.6]
  wire  loadRequest_4; // @[LoadQueue.scala 229:71:@40764.4]
  wire [15:0] _T_90467; // @[Mux.scala 31:69:@39170.4]
  wire  _T_92504; // @[LoadQueue.scala 229:41:@40680.4]
  wire  _T_92505; // @[LoadQueue.scala 229:38:@40681.4]
  wire  _T_92507; // @[LoadQueue.scala 230:12:@40683.6]
  reg  prevPriorityRequest_3; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_751;
  wire  _T_92509; // @[LoadQueue.scala 230:46:@40684.6]
  wire  _T_92510; // @[LoadQueue.scala 230:43:@40685.6]
  wire  _T_92512; // @[LoadQueue.scala 230:84:@40686.6]
  wire  _T_92513; // @[LoadQueue.scala 230:81:@40687.6]
  wire  _T_92516; // @[LoadQueue.scala 233:86:@40690.8]
  wire  _T_92517; // @[LoadQueue.scala 233:86:@40691.8]
  wire  _T_92518; // @[LoadQueue.scala 233:86:@40692.8]
  wire  _T_92519; // @[LoadQueue.scala 233:86:@40693.8]
  wire  _T_92520; // @[LoadQueue.scala 233:86:@40694.8]
  wire  _T_92521; // @[LoadQueue.scala 233:86:@40695.8]
  wire  _T_92522; // @[LoadQueue.scala 233:86:@40696.8]
  wire  _T_92523; // @[LoadQueue.scala 233:86:@40697.8]
  wire  _T_92524; // @[LoadQueue.scala 233:86:@40698.8]
  wire  _T_92525; // @[LoadQueue.scala 233:86:@40699.8]
  wire  _T_92526; // @[LoadQueue.scala 233:86:@40700.8]
  wire  _T_92527; // @[LoadQueue.scala 233:86:@40701.8]
  wire  _T_92528; // @[LoadQueue.scala 233:86:@40702.8]
  wire  _T_92529; // @[LoadQueue.scala 233:86:@40703.8]
  wire  _T_92530; // @[LoadQueue.scala 233:86:@40704.8]
  wire  _T_92532; // @[LoadQueue.scala 233:38:@40705.8]
  wire  _T_92551; // @[LoadQueue.scala 234:11:@40722.8]
  wire  _T_92552; // @[LoadQueue.scala 233:103:@40723.8]
  wire  _GEN_1980; // @[LoadQueue.scala 230:110:@40688.6]
  wire  loadRequest_3; // @[LoadQueue.scala 229:71:@40682.4]
  wire [15:0] _T_90468; // @[Mux.scala 31:69:@39171.4]
  wire  _T_92420; // @[LoadQueue.scala 229:41:@40598.4]
  wire  _T_92421; // @[LoadQueue.scala 229:38:@40599.4]
  wire  _T_92423; // @[LoadQueue.scala 230:12:@40601.6]
  reg  prevPriorityRequest_2; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_752;
  wire  _T_92425; // @[LoadQueue.scala 230:46:@40602.6]
  wire  _T_92426; // @[LoadQueue.scala 230:43:@40603.6]
  wire  _T_92428; // @[LoadQueue.scala 230:84:@40604.6]
  wire  _T_92429; // @[LoadQueue.scala 230:81:@40605.6]
  wire  _T_92432; // @[LoadQueue.scala 233:86:@40608.8]
  wire  _T_92433; // @[LoadQueue.scala 233:86:@40609.8]
  wire  _T_92434; // @[LoadQueue.scala 233:86:@40610.8]
  wire  _T_92435; // @[LoadQueue.scala 233:86:@40611.8]
  wire  _T_92436; // @[LoadQueue.scala 233:86:@40612.8]
  wire  _T_92437; // @[LoadQueue.scala 233:86:@40613.8]
  wire  _T_92438; // @[LoadQueue.scala 233:86:@40614.8]
  wire  _T_92439; // @[LoadQueue.scala 233:86:@40615.8]
  wire  _T_92440; // @[LoadQueue.scala 233:86:@40616.8]
  wire  _T_92441; // @[LoadQueue.scala 233:86:@40617.8]
  wire  _T_92442; // @[LoadQueue.scala 233:86:@40618.8]
  wire  _T_92443; // @[LoadQueue.scala 233:86:@40619.8]
  wire  _T_92444; // @[LoadQueue.scala 233:86:@40620.8]
  wire  _T_92445; // @[LoadQueue.scala 233:86:@40621.8]
  wire  _T_92446; // @[LoadQueue.scala 233:86:@40622.8]
  wire  _T_92448; // @[LoadQueue.scala 233:38:@40623.8]
  wire  _T_92467; // @[LoadQueue.scala 234:11:@40640.8]
  wire  _T_92468; // @[LoadQueue.scala 233:103:@40641.8]
  wire  _GEN_1976; // @[LoadQueue.scala 230:110:@40606.6]
  wire  loadRequest_2; // @[LoadQueue.scala 229:71:@40600.4]
  wire [15:0] _T_90469; // @[Mux.scala 31:69:@39172.4]
  wire  _T_92336; // @[LoadQueue.scala 229:41:@40516.4]
  wire  _T_92337; // @[LoadQueue.scala 229:38:@40517.4]
  wire  _T_92339; // @[LoadQueue.scala 230:12:@40519.6]
  reg  prevPriorityRequest_1; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_753;
  wire  _T_92341; // @[LoadQueue.scala 230:46:@40520.6]
  wire  _T_92342; // @[LoadQueue.scala 230:43:@40521.6]
  wire  _T_92344; // @[LoadQueue.scala 230:84:@40522.6]
  wire  _T_92345; // @[LoadQueue.scala 230:81:@40523.6]
  wire  _T_92348; // @[LoadQueue.scala 233:86:@40526.8]
  wire  _T_92349; // @[LoadQueue.scala 233:86:@40527.8]
  wire  _T_92350; // @[LoadQueue.scala 233:86:@40528.8]
  wire  _T_92351; // @[LoadQueue.scala 233:86:@40529.8]
  wire  _T_92352; // @[LoadQueue.scala 233:86:@40530.8]
  wire  _T_92353; // @[LoadQueue.scala 233:86:@40531.8]
  wire  _T_92354; // @[LoadQueue.scala 233:86:@40532.8]
  wire  _T_92355; // @[LoadQueue.scala 233:86:@40533.8]
  wire  _T_92356; // @[LoadQueue.scala 233:86:@40534.8]
  wire  _T_92357; // @[LoadQueue.scala 233:86:@40535.8]
  wire  _T_92358; // @[LoadQueue.scala 233:86:@40536.8]
  wire  _T_92359; // @[LoadQueue.scala 233:86:@40537.8]
  wire  _T_92360; // @[LoadQueue.scala 233:86:@40538.8]
  wire  _T_92361; // @[LoadQueue.scala 233:86:@40539.8]
  wire  _T_92362; // @[LoadQueue.scala 233:86:@40540.8]
  wire  _T_92364; // @[LoadQueue.scala 233:38:@40541.8]
  wire  _T_92383; // @[LoadQueue.scala 234:11:@40558.8]
  wire  _T_92384; // @[LoadQueue.scala 233:103:@40559.8]
  wire  _GEN_1972; // @[LoadQueue.scala 230:110:@40524.6]
  wire  loadRequest_1; // @[LoadQueue.scala 229:71:@40518.4]
  wire [15:0] _T_90470; // @[Mux.scala 31:69:@39173.4]
  wire  _T_92252; // @[LoadQueue.scala 229:41:@40434.4]
  wire  _T_92253; // @[LoadQueue.scala 229:38:@40435.4]
  wire  _T_92255; // @[LoadQueue.scala 230:12:@40437.6]
  reg  prevPriorityRequest_0; // @[LoadQueue.scala 207:36:@40266.4]
  reg [31:0] _RAND_754;
  wire  _T_92257; // @[LoadQueue.scala 230:46:@40438.6]
  wire  _T_92258; // @[LoadQueue.scala 230:43:@40439.6]
  wire  _T_92260; // @[LoadQueue.scala 230:84:@40440.6]
  wire  _T_92261; // @[LoadQueue.scala 230:81:@40441.6]
  wire  _T_92264; // @[LoadQueue.scala 233:86:@40444.8]
  wire  _T_92265; // @[LoadQueue.scala 233:86:@40445.8]
  wire  _T_92266; // @[LoadQueue.scala 233:86:@40446.8]
  wire  _T_92267; // @[LoadQueue.scala 233:86:@40447.8]
  wire  _T_92268; // @[LoadQueue.scala 233:86:@40448.8]
  wire  _T_92269; // @[LoadQueue.scala 233:86:@40449.8]
  wire  _T_92270; // @[LoadQueue.scala 233:86:@40450.8]
  wire  _T_92271; // @[LoadQueue.scala 233:86:@40451.8]
  wire  _T_92272; // @[LoadQueue.scala 233:86:@40452.8]
  wire  _T_92273; // @[LoadQueue.scala 233:86:@40453.8]
  wire  _T_92274; // @[LoadQueue.scala 233:86:@40454.8]
  wire  _T_92275; // @[LoadQueue.scala 233:86:@40455.8]
  wire  _T_92276; // @[LoadQueue.scala 233:86:@40456.8]
  wire  _T_92277; // @[LoadQueue.scala 233:86:@40457.8]
  wire  _T_92278; // @[LoadQueue.scala 233:86:@40458.8]
  wire  _T_92280; // @[LoadQueue.scala 233:38:@40459.8]
  wire  _T_92299; // @[LoadQueue.scala 234:11:@40476.8]
  wire  _T_92300; // @[LoadQueue.scala 233:103:@40477.8]
  wire  _GEN_1968; // @[LoadQueue.scala 230:110:@40442.6]
  wire  loadRequest_0; // @[LoadQueue.scala 229:71:@40436.4]
  wire [15:0] _T_90471; // @[Mux.scala 31:69:@39174.4]
  wire  _T_90472; // @[OneHot.scala 66:30:@39175.4]
  wire  _T_90473; // @[OneHot.scala 66:30:@39176.4]
  wire  _T_90474; // @[OneHot.scala 66:30:@39177.4]
  wire  _T_90475; // @[OneHot.scala 66:30:@39178.4]
  wire  _T_90476; // @[OneHot.scala 66:30:@39179.4]
  wire  _T_90477; // @[OneHot.scala 66:30:@39180.4]
  wire  _T_90478; // @[OneHot.scala 66:30:@39181.4]
  wire  _T_90479; // @[OneHot.scala 66:30:@39182.4]
  wire  _T_90480; // @[OneHot.scala 66:30:@39183.4]
  wire  _T_90481; // @[OneHot.scala 66:30:@39184.4]
  wire  _T_90482; // @[OneHot.scala 66:30:@39185.4]
  wire  _T_90483; // @[OneHot.scala 66:30:@39186.4]
  wire  _T_90484; // @[OneHot.scala 66:30:@39187.4]
  wire  _T_90485; // @[OneHot.scala 66:30:@39188.4]
  wire  _T_90486; // @[OneHot.scala 66:30:@39189.4]
  wire  _T_90487; // @[OneHot.scala 66:30:@39190.4]
  wire [15:0] _T_90528; // @[Mux.scala 31:69:@39208.4]
  wire [15:0] _T_90529; // @[Mux.scala 31:69:@39209.4]
  wire [15:0] _T_90530; // @[Mux.scala 31:69:@39210.4]
  wire [15:0] _T_90531; // @[Mux.scala 31:69:@39211.4]
  wire [15:0] _T_90532; // @[Mux.scala 31:69:@39212.4]
  wire [15:0] _T_90533; // @[Mux.scala 31:69:@39213.4]
  wire [15:0] _T_90534; // @[Mux.scala 31:69:@39214.4]
  wire [15:0] _T_90535; // @[Mux.scala 31:69:@39215.4]
  wire [15:0] _T_90536; // @[Mux.scala 31:69:@39216.4]
  wire [15:0] _T_90537; // @[Mux.scala 31:69:@39217.4]
  wire [15:0] _T_90538; // @[Mux.scala 31:69:@39218.4]
  wire [15:0] _T_90539; // @[Mux.scala 31:69:@39219.4]
  wire [15:0] _T_90540; // @[Mux.scala 31:69:@39220.4]
  wire [15:0] _T_90541; // @[Mux.scala 31:69:@39221.4]
  wire [15:0] _T_90542; // @[Mux.scala 31:69:@39222.4]
  wire [15:0] _T_90543; // @[Mux.scala 31:69:@39223.4]
  wire  _T_90544; // @[OneHot.scala 66:30:@39224.4]
  wire  _T_90545; // @[OneHot.scala 66:30:@39225.4]
  wire  _T_90546; // @[OneHot.scala 66:30:@39226.4]
  wire  _T_90547; // @[OneHot.scala 66:30:@39227.4]
  wire  _T_90548; // @[OneHot.scala 66:30:@39228.4]
  wire  _T_90549; // @[OneHot.scala 66:30:@39229.4]
  wire  _T_90550; // @[OneHot.scala 66:30:@39230.4]
  wire  _T_90551; // @[OneHot.scala 66:30:@39231.4]
  wire  _T_90552; // @[OneHot.scala 66:30:@39232.4]
  wire  _T_90553; // @[OneHot.scala 66:30:@39233.4]
  wire  _T_90554; // @[OneHot.scala 66:30:@39234.4]
  wire  _T_90555; // @[OneHot.scala 66:30:@39235.4]
  wire  _T_90556; // @[OneHot.scala 66:30:@39236.4]
  wire  _T_90557; // @[OneHot.scala 66:30:@39237.4]
  wire  _T_90558; // @[OneHot.scala 66:30:@39238.4]
  wire  _T_90559; // @[OneHot.scala 66:30:@39239.4]
  wire [15:0] _T_90600; // @[Mux.scala 31:69:@39257.4]
  wire [15:0] _T_90601; // @[Mux.scala 31:69:@39258.4]
  wire [15:0] _T_90602; // @[Mux.scala 31:69:@39259.4]
  wire [15:0] _T_90603; // @[Mux.scala 31:69:@39260.4]
  wire [15:0] _T_90604; // @[Mux.scala 31:69:@39261.4]
  wire [15:0] _T_90605; // @[Mux.scala 31:69:@39262.4]
  wire [15:0] _T_90606; // @[Mux.scala 31:69:@39263.4]
  wire [15:0] _T_90607; // @[Mux.scala 31:69:@39264.4]
  wire [15:0] _T_90608; // @[Mux.scala 31:69:@39265.4]
  wire [15:0] _T_90609; // @[Mux.scala 31:69:@39266.4]
  wire [15:0] _T_90610; // @[Mux.scala 31:69:@39267.4]
  wire [15:0] _T_90611; // @[Mux.scala 31:69:@39268.4]
  wire [15:0] _T_90612; // @[Mux.scala 31:69:@39269.4]
  wire [15:0] _T_90613; // @[Mux.scala 31:69:@39270.4]
  wire [15:0] _T_90614; // @[Mux.scala 31:69:@39271.4]
  wire [15:0] _T_90615; // @[Mux.scala 31:69:@39272.4]
  wire  _T_90616; // @[OneHot.scala 66:30:@39273.4]
  wire  _T_90617; // @[OneHot.scala 66:30:@39274.4]
  wire  _T_90618; // @[OneHot.scala 66:30:@39275.4]
  wire  _T_90619; // @[OneHot.scala 66:30:@39276.4]
  wire  _T_90620; // @[OneHot.scala 66:30:@39277.4]
  wire  _T_90621; // @[OneHot.scala 66:30:@39278.4]
  wire  _T_90622; // @[OneHot.scala 66:30:@39279.4]
  wire  _T_90623; // @[OneHot.scala 66:30:@39280.4]
  wire  _T_90624; // @[OneHot.scala 66:30:@39281.4]
  wire  _T_90625; // @[OneHot.scala 66:30:@39282.4]
  wire  _T_90626; // @[OneHot.scala 66:30:@39283.4]
  wire  _T_90627; // @[OneHot.scala 66:30:@39284.4]
  wire  _T_90628; // @[OneHot.scala 66:30:@39285.4]
  wire  _T_90629; // @[OneHot.scala 66:30:@39286.4]
  wire  _T_90630; // @[OneHot.scala 66:30:@39287.4]
  wire  _T_90631; // @[OneHot.scala 66:30:@39288.4]
  wire [15:0] _T_90672; // @[Mux.scala 31:69:@39306.4]
  wire [15:0] _T_90673; // @[Mux.scala 31:69:@39307.4]
  wire [15:0] _T_90674; // @[Mux.scala 31:69:@39308.4]
  wire [15:0] _T_90675; // @[Mux.scala 31:69:@39309.4]
  wire [15:0] _T_90676; // @[Mux.scala 31:69:@39310.4]
  wire [15:0] _T_90677; // @[Mux.scala 31:69:@39311.4]
  wire [15:0] _T_90678; // @[Mux.scala 31:69:@39312.4]
  wire [15:0] _T_90679; // @[Mux.scala 31:69:@39313.4]
  wire [15:0] _T_90680; // @[Mux.scala 31:69:@39314.4]
  wire [15:0] _T_90681; // @[Mux.scala 31:69:@39315.4]
  wire [15:0] _T_90682; // @[Mux.scala 31:69:@39316.4]
  wire [15:0] _T_90683; // @[Mux.scala 31:69:@39317.4]
  wire [15:0] _T_90684; // @[Mux.scala 31:69:@39318.4]
  wire [15:0] _T_90685; // @[Mux.scala 31:69:@39319.4]
  wire [15:0] _T_90686; // @[Mux.scala 31:69:@39320.4]
  wire [15:0] _T_90687; // @[Mux.scala 31:69:@39321.4]
  wire  _T_90688; // @[OneHot.scala 66:30:@39322.4]
  wire  _T_90689; // @[OneHot.scala 66:30:@39323.4]
  wire  _T_90690; // @[OneHot.scala 66:30:@39324.4]
  wire  _T_90691; // @[OneHot.scala 66:30:@39325.4]
  wire  _T_90692; // @[OneHot.scala 66:30:@39326.4]
  wire  _T_90693; // @[OneHot.scala 66:30:@39327.4]
  wire  _T_90694; // @[OneHot.scala 66:30:@39328.4]
  wire  _T_90695; // @[OneHot.scala 66:30:@39329.4]
  wire  _T_90696; // @[OneHot.scala 66:30:@39330.4]
  wire  _T_90697; // @[OneHot.scala 66:30:@39331.4]
  wire  _T_90698; // @[OneHot.scala 66:30:@39332.4]
  wire  _T_90699; // @[OneHot.scala 66:30:@39333.4]
  wire  _T_90700; // @[OneHot.scala 66:30:@39334.4]
  wire  _T_90701; // @[OneHot.scala 66:30:@39335.4]
  wire  _T_90702; // @[OneHot.scala 66:30:@39336.4]
  wire  _T_90703; // @[OneHot.scala 66:30:@39337.4]
  wire [15:0] _T_90744; // @[Mux.scala 31:69:@39355.4]
  wire [15:0] _T_90745; // @[Mux.scala 31:69:@39356.4]
  wire [15:0] _T_90746; // @[Mux.scala 31:69:@39357.4]
  wire [15:0] _T_90747; // @[Mux.scala 31:69:@39358.4]
  wire [15:0] _T_90748; // @[Mux.scala 31:69:@39359.4]
  wire [15:0] _T_90749; // @[Mux.scala 31:69:@39360.4]
  wire [15:0] _T_90750; // @[Mux.scala 31:69:@39361.4]
  wire [15:0] _T_90751; // @[Mux.scala 31:69:@39362.4]
  wire [15:0] _T_90752; // @[Mux.scala 31:69:@39363.4]
  wire [15:0] _T_90753; // @[Mux.scala 31:69:@39364.4]
  wire [15:0] _T_90754; // @[Mux.scala 31:69:@39365.4]
  wire [15:0] _T_90755; // @[Mux.scala 31:69:@39366.4]
  wire [15:0] _T_90756; // @[Mux.scala 31:69:@39367.4]
  wire [15:0] _T_90757; // @[Mux.scala 31:69:@39368.4]
  wire [15:0] _T_90758; // @[Mux.scala 31:69:@39369.4]
  wire [15:0] _T_90759; // @[Mux.scala 31:69:@39370.4]
  wire  _T_90760; // @[OneHot.scala 66:30:@39371.4]
  wire  _T_90761; // @[OneHot.scala 66:30:@39372.4]
  wire  _T_90762; // @[OneHot.scala 66:30:@39373.4]
  wire  _T_90763; // @[OneHot.scala 66:30:@39374.4]
  wire  _T_90764; // @[OneHot.scala 66:30:@39375.4]
  wire  _T_90765; // @[OneHot.scala 66:30:@39376.4]
  wire  _T_90766; // @[OneHot.scala 66:30:@39377.4]
  wire  _T_90767; // @[OneHot.scala 66:30:@39378.4]
  wire  _T_90768; // @[OneHot.scala 66:30:@39379.4]
  wire  _T_90769; // @[OneHot.scala 66:30:@39380.4]
  wire  _T_90770; // @[OneHot.scala 66:30:@39381.4]
  wire  _T_90771; // @[OneHot.scala 66:30:@39382.4]
  wire  _T_90772; // @[OneHot.scala 66:30:@39383.4]
  wire  _T_90773; // @[OneHot.scala 66:30:@39384.4]
  wire  _T_90774; // @[OneHot.scala 66:30:@39385.4]
  wire  _T_90775; // @[OneHot.scala 66:30:@39386.4]
  wire [15:0] _T_90816; // @[Mux.scala 31:69:@39404.4]
  wire [15:0] _T_90817; // @[Mux.scala 31:69:@39405.4]
  wire [15:0] _T_90818; // @[Mux.scala 31:69:@39406.4]
  wire [15:0] _T_90819; // @[Mux.scala 31:69:@39407.4]
  wire [15:0] _T_90820; // @[Mux.scala 31:69:@39408.4]
  wire [15:0] _T_90821; // @[Mux.scala 31:69:@39409.4]
  wire [15:0] _T_90822; // @[Mux.scala 31:69:@39410.4]
  wire [15:0] _T_90823; // @[Mux.scala 31:69:@39411.4]
  wire [15:0] _T_90824; // @[Mux.scala 31:69:@39412.4]
  wire [15:0] _T_90825; // @[Mux.scala 31:69:@39413.4]
  wire [15:0] _T_90826; // @[Mux.scala 31:69:@39414.4]
  wire [15:0] _T_90827; // @[Mux.scala 31:69:@39415.4]
  wire [15:0] _T_90828; // @[Mux.scala 31:69:@39416.4]
  wire [15:0] _T_90829; // @[Mux.scala 31:69:@39417.4]
  wire [15:0] _T_90830; // @[Mux.scala 31:69:@39418.4]
  wire [15:0] _T_90831; // @[Mux.scala 31:69:@39419.4]
  wire  _T_90832; // @[OneHot.scala 66:30:@39420.4]
  wire  _T_90833; // @[OneHot.scala 66:30:@39421.4]
  wire  _T_90834; // @[OneHot.scala 66:30:@39422.4]
  wire  _T_90835; // @[OneHot.scala 66:30:@39423.4]
  wire  _T_90836; // @[OneHot.scala 66:30:@39424.4]
  wire  _T_90837; // @[OneHot.scala 66:30:@39425.4]
  wire  _T_90838; // @[OneHot.scala 66:30:@39426.4]
  wire  _T_90839; // @[OneHot.scala 66:30:@39427.4]
  wire  _T_90840; // @[OneHot.scala 66:30:@39428.4]
  wire  _T_90841; // @[OneHot.scala 66:30:@39429.4]
  wire  _T_90842; // @[OneHot.scala 66:30:@39430.4]
  wire  _T_90843; // @[OneHot.scala 66:30:@39431.4]
  wire  _T_90844; // @[OneHot.scala 66:30:@39432.4]
  wire  _T_90845; // @[OneHot.scala 66:30:@39433.4]
  wire  _T_90846; // @[OneHot.scala 66:30:@39434.4]
  wire  _T_90847; // @[OneHot.scala 66:30:@39435.4]
  wire [15:0] _T_90888; // @[Mux.scala 31:69:@39453.4]
  wire [15:0] _T_90889; // @[Mux.scala 31:69:@39454.4]
  wire [15:0] _T_90890; // @[Mux.scala 31:69:@39455.4]
  wire [15:0] _T_90891; // @[Mux.scala 31:69:@39456.4]
  wire [15:0] _T_90892; // @[Mux.scala 31:69:@39457.4]
  wire [15:0] _T_90893; // @[Mux.scala 31:69:@39458.4]
  wire [15:0] _T_90894; // @[Mux.scala 31:69:@39459.4]
  wire [15:0] _T_90895; // @[Mux.scala 31:69:@39460.4]
  wire [15:0] _T_90896; // @[Mux.scala 31:69:@39461.4]
  wire [15:0] _T_90897; // @[Mux.scala 31:69:@39462.4]
  wire [15:0] _T_90898; // @[Mux.scala 31:69:@39463.4]
  wire [15:0] _T_90899; // @[Mux.scala 31:69:@39464.4]
  wire [15:0] _T_90900; // @[Mux.scala 31:69:@39465.4]
  wire [15:0] _T_90901; // @[Mux.scala 31:69:@39466.4]
  wire [15:0] _T_90902; // @[Mux.scala 31:69:@39467.4]
  wire [15:0] _T_90903; // @[Mux.scala 31:69:@39468.4]
  wire  _T_90904; // @[OneHot.scala 66:30:@39469.4]
  wire  _T_90905; // @[OneHot.scala 66:30:@39470.4]
  wire  _T_90906; // @[OneHot.scala 66:30:@39471.4]
  wire  _T_90907; // @[OneHot.scala 66:30:@39472.4]
  wire  _T_90908; // @[OneHot.scala 66:30:@39473.4]
  wire  _T_90909; // @[OneHot.scala 66:30:@39474.4]
  wire  _T_90910; // @[OneHot.scala 66:30:@39475.4]
  wire  _T_90911; // @[OneHot.scala 66:30:@39476.4]
  wire  _T_90912; // @[OneHot.scala 66:30:@39477.4]
  wire  _T_90913; // @[OneHot.scala 66:30:@39478.4]
  wire  _T_90914; // @[OneHot.scala 66:30:@39479.4]
  wire  _T_90915; // @[OneHot.scala 66:30:@39480.4]
  wire  _T_90916; // @[OneHot.scala 66:30:@39481.4]
  wire  _T_90917; // @[OneHot.scala 66:30:@39482.4]
  wire  _T_90918; // @[OneHot.scala 66:30:@39483.4]
  wire  _T_90919; // @[OneHot.scala 66:30:@39484.4]
  wire [15:0] _T_90960; // @[Mux.scala 31:69:@39502.4]
  wire [15:0] _T_90961; // @[Mux.scala 31:69:@39503.4]
  wire [15:0] _T_90962; // @[Mux.scala 31:69:@39504.4]
  wire [15:0] _T_90963; // @[Mux.scala 31:69:@39505.4]
  wire [15:0] _T_90964; // @[Mux.scala 31:69:@39506.4]
  wire [15:0] _T_90965; // @[Mux.scala 31:69:@39507.4]
  wire [15:0] _T_90966; // @[Mux.scala 31:69:@39508.4]
  wire [15:0] _T_90967; // @[Mux.scala 31:69:@39509.4]
  wire [15:0] _T_90968; // @[Mux.scala 31:69:@39510.4]
  wire [15:0] _T_90969; // @[Mux.scala 31:69:@39511.4]
  wire [15:0] _T_90970; // @[Mux.scala 31:69:@39512.4]
  wire [15:0] _T_90971; // @[Mux.scala 31:69:@39513.4]
  wire [15:0] _T_90972; // @[Mux.scala 31:69:@39514.4]
  wire [15:0] _T_90973; // @[Mux.scala 31:69:@39515.4]
  wire [15:0] _T_90974; // @[Mux.scala 31:69:@39516.4]
  wire [15:0] _T_90975; // @[Mux.scala 31:69:@39517.4]
  wire  _T_90976; // @[OneHot.scala 66:30:@39518.4]
  wire  _T_90977; // @[OneHot.scala 66:30:@39519.4]
  wire  _T_90978; // @[OneHot.scala 66:30:@39520.4]
  wire  _T_90979; // @[OneHot.scala 66:30:@39521.4]
  wire  _T_90980; // @[OneHot.scala 66:30:@39522.4]
  wire  _T_90981; // @[OneHot.scala 66:30:@39523.4]
  wire  _T_90982; // @[OneHot.scala 66:30:@39524.4]
  wire  _T_90983; // @[OneHot.scala 66:30:@39525.4]
  wire  _T_90984; // @[OneHot.scala 66:30:@39526.4]
  wire  _T_90985; // @[OneHot.scala 66:30:@39527.4]
  wire  _T_90986; // @[OneHot.scala 66:30:@39528.4]
  wire  _T_90987; // @[OneHot.scala 66:30:@39529.4]
  wire  _T_90988; // @[OneHot.scala 66:30:@39530.4]
  wire  _T_90989; // @[OneHot.scala 66:30:@39531.4]
  wire  _T_90990; // @[OneHot.scala 66:30:@39532.4]
  wire  _T_90991; // @[OneHot.scala 66:30:@39533.4]
  wire [15:0] _T_91032; // @[Mux.scala 31:69:@39551.4]
  wire [15:0] _T_91033; // @[Mux.scala 31:69:@39552.4]
  wire [15:0] _T_91034; // @[Mux.scala 31:69:@39553.4]
  wire [15:0] _T_91035; // @[Mux.scala 31:69:@39554.4]
  wire [15:0] _T_91036; // @[Mux.scala 31:69:@39555.4]
  wire [15:0] _T_91037; // @[Mux.scala 31:69:@39556.4]
  wire [15:0] _T_91038; // @[Mux.scala 31:69:@39557.4]
  wire [15:0] _T_91039; // @[Mux.scala 31:69:@39558.4]
  wire [15:0] _T_91040; // @[Mux.scala 31:69:@39559.4]
  wire [15:0] _T_91041; // @[Mux.scala 31:69:@39560.4]
  wire [15:0] _T_91042; // @[Mux.scala 31:69:@39561.4]
  wire [15:0] _T_91043; // @[Mux.scala 31:69:@39562.4]
  wire [15:0] _T_91044; // @[Mux.scala 31:69:@39563.4]
  wire [15:0] _T_91045; // @[Mux.scala 31:69:@39564.4]
  wire [15:0] _T_91046; // @[Mux.scala 31:69:@39565.4]
  wire [15:0] _T_91047; // @[Mux.scala 31:69:@39566.4]
  wire  _T_91048; // @[OneHot.scala 66:30:@39567.4]
  wire  _T_91049; // @[OneHot.scala 66:30:@39568.4]
  wire  _T_91050; // @[OneHot.scala 66:30:@39569.4]
  wire  _T_91051; // @[OneHot.scala 66:30:@39570.4]
  wire  _T_91052; // @[OneHot.scala 66:30:@39571.4]
  wire  _T_91053; // @[OneHot.scala 66:30:@39572.4]
  wire  _T_91054; // @[OneHot.scala 66:30:@39573.4]
  wire  _T_91055; // @[OneHot.scala 66:30:@39574.4]
  wire  _T_91056; // @[OneHot.scala 66:30:@39575.4]
  wire  _T_91057; // @[OneHot.scala 66:30:@39576.4]
  wire  _T_91058; // @[OneHot.scala 66:30:@39577.4]
  wire  _T_91059; // @[OneHot.scala 66:30:@39578.4]
  wire  _T_91060; // @[OneHot.scala 66:30:@39579.4]
  wire  _T_91061; // @[OneHot.scala 66:30:@39580.4]
  wire  _T_91062; // @[OneHot.scala 66:30:@39581.4]
  wire  _T_91063; // @[OneHot.scala 66:30:@39582.4]
  wire [15:0] _T_91104; // @[Mux.scala 31:69:@39600.4]
  wire [15:0] _T_91105; // @[Mux.scala 31:69:@39601.4]
  wire [15:0] _T_91106; // @[Mux.scala 31:69:@39602.4]
  wire [15:0] _T_91107; // @[Mux.scala 31:69:@39603.4]
  wire [15:0] _T_91108; // @[Mux.scala 31:69:@39604.4]
  wire [15:0] _T_91109; // @[Mux.scala 31:69:@39605.4]
  wire [15:0] _T_91110; // @[Mux.scala 31:69:@39606.4]
  wire [15:0] _T_91111; // @[Mux.scala 31:69:@39607.4]
  wire [15:0] _T_91112; // @[Mux.scala 31:69:@39608.4]
  wire [15:0] _T_91113; // @[Mux.scala 31:69:@39609.4]
  wire [15:0] _T_91114; // @[Mux.scala 31:69:@39610.4]
  wire [15:0] _T_91115; // @[Mux.scala 31:69:@39611.4]
  wire [15:0] _T_91116; // @[Mux.scala 31:69:@39612.4]
  wire [15:0] _T_91117; // @[Mux.scala 31:69:@39613.4]
  wire [15:0] _T_91118; // @[Mux.scala 31:69:@39614.4]
  wire [15:0] _T_91119; // @[Mux.scala 31:69:@39615.4]
  wire  _T_91120; // @[OneHot.scala 66:30:@39616.4]
  wire  _T_91121; // @[OneHot.scala 66:30:@39617.4]
  wire  _T_91122; // @[OneHot.scala 66:30:@39618.4]
  wire  _T_91123; // @[OneHot.scala 66:30:@39619.4]
  wire  _T_91124; // @[OneHot.scala 66:30:@39620.4]
  wire  _T_91125; // @[OneHot.scala 66:30:@39621.4]
  wire  _T_91126; // @[OneHot.scala 66:30:@39622.4]
  wire  _T_91127; // @[OneHot.scala 66:30:@39623.4]
  wire  _T_91128; // @[OneHot.scala 66:30:@39624.4]
  wire  _T_91129; // @[OneHot.scala 66:30:@39625.4]
  wire  _T_91130; // @[OneHot.scala 66:30:@39626.4]
  wire  _T_91131; // @[OneHot.scala 66:30:@39627.4]
  wire  _T_91132; // @[OneHot.scala 66:30:@39628.4]
  wire  _T_91133; // @[OneHot.scala 66:30:@39629.4]
  wire  _T_91134; // @[OneHot.scala 66:30:@39630.4]
  wire  _T_91135; // @[OneHot.scala 66:30:@39631.4]
  wire [15:0] _T_91176; // @[Mux.scala 31:69:@39649.4]
  wire [15:0] _T_91177; // @[Mux.scala 31:69:@39650.4]
  wire [15:0] _T_91178; // @[Mux.scala 31:69:@39651.4]
  wire [15:0] _T_91179; // @[Mux.scala 31:69:@39652.4]
  wire [15:0] _T_91180; // @[Mux.scala 31:69:@39653.4]
  wire [15:0] _T_91181; // @[Mux.scala 31:69:@39654.4]
  wire [15:0] _T_91182; // @[Mux.scala 31:69:@39655.4]
  wire [15:0] _T_91183; // @[Mux.scala 31:69:@39656.4]
  wire [15:0] _T_91184; // @[Mux.scala 31:69:@39657.4]
  wire [15:0] _T_91185; // @[Mux.scala 31:69:@39658.4]
  wire [15:0] _T_91186; // @[Mux.scala 31:69:@39659.4]
  wire [15:0] _T_91187; // @[Mux.scala 31:69:@39660.4]
  wire [15:0] _T_91188; // @[Mux.scala 31:69:@39661.4]
  wire [15:0] _T_91189; // @[Mux.scala 31:69:@39662.4]
  wire [15:0] _T_91190; // @[Mux.scala 31:69:@39663.4]
  wire [15:0] _T_91191; // @[Mux.scala 31:69:@39664.4]
  wire  _T_91192; // @[OneHot.scala 66:30:@39665.4]
  wire  _T_91193; // @[OneHot.scala 66:30:@39666.4]
  wire  _T_91194; // @[OneHot.scala 66:30:@39667.4]
  wire  _T_91195; // @[OneHot.scala 66:30:@39668.4]
  wire  _T_91196; // @[OneHot.scala 66:30:@39669.4]
  wire  _T_91197; // @[OneHot.scala 66:30:@39670.4]
  wire  _T_91198; // @[OneHot.scala 66:30:@39671.4]
  wire  _T_91199; // @[OneHot.scala 66:30:@39672.4]
  wire  _T_91200; // @[OneHot.scala 66:30:@39673.4]
  wire  _T_91201; // @[OneHot.scala 66:30:@39674.4]
  wire  _T_91202; // @[OneHot.scala 66:30:@39675.4]
  wire  _T_91203; // @[OneHot.scala 66:30:@39676.4]
  wire  _T_91204; // @[OneHot.scala 66:30:@39677.4]
  wire  _T_91205; // @[OneHot.scala 66:30:@39678.4]
  wire  _T_91206; // @[OneHot.scala 66:30:@39679.4]
  wire  _T_91207; // @[OneHot.scala 66:30:@39680.4]
  wire [15:0] _T_91248; // @[Mux.scala 31:69:@39698.4]
  wire [15:0] _T_91249; // @[Mux.scala 31:69:@39699.4]
  wire [15:0] _T_91250; // @[Mux.scala 31:69:@39700.4]
  wire [15:0] _T_91251; // @[Mux.scala 31:69:@39701.4]
  wire [15:0] _T_91252; // @[Mux.scala 31:69:@39702.4]
  wire [15:0] _T_91253; // @[Mux.scala 31:69:@39703.4]
  wire [15:0] _T_91254; // @[Mux.scala 31:69:@39704.4]
  wire [15:0] _T_91255; // @[Mux.scala 31:69:@39705.4]
  wire [15:0] _T_91256; // @[Mux.scala 31:69:@39706.4]
  wire [15:0] _T_91257; // @[Mux.scala 31:69:@39707.4]
  wire [15:0] _T_91258; // @[Mux.scala 31:69:@39708.4]
  wire [15:0] _T_91259; // @[Mux.scala 31:69:@39709.4]
  wire [15:0] _T_91260; // @[Mux.scala 31:69:@39710.4]
  wire [15:0] _T_91261; // @[Mux.scala 31:69:@39711.4]
  wire [15:0] _T_91262; // @[Mux.scala 31:69:@39712.4]
  wire [15:0] _T_91263; // @[Mux.scala 31:69:@39713.4]
  wire  _T_91264; // @[OneHot.scala 66:30:@39714.4]
  wire  _T_91265; // @[OneHot.scala 66:30:@39715.4]
  wire  _T_91266; // @[OneHot.scala 66:30:@39716.4]
  wire  _T_91267; // @[OneHot.scala 66:30:@39717.4]
  wire  _T_91268; // @[OneHot.scala 66:30:@39718.4]
  wire  _T_91269; // @[OneHot.scala 66:30:@39719.4]
  wire  _T_91270; // @[OneHot.scala 66:30:@39720.4]
  wire  _T_91271; // @[OneHot.scala 66:30:@39721.4]
  wire  _T_91272; // @[OneHot.scala 66:30:@39722.4]
  wire  _T_91273; // @[OneHot.scala 66:30:@39723.4]
  wire  _T_91274; // @[OneHot.scala 66:30:@39724.4]
  wire  _T_91275; // @[OneHot.scala 66:30:@39725.4]
  wire  _T_91276; // @[OneHot.scala 66:30:@39726.4]
  wire  _T_91277; // @[OneHot.scala 66:30:@39727.4]
  wire  _T_91278; // @[OneHot.scala 66:30:@39728.4]
  wire  _T_91279; // @[OneHot.scala 66:30:@39729.4]
  wire [15:0] _T_91320; // @[Mux.scala 31:69:@39747.4]
  wire [15:0] _T_91321; // @[Mux.scala 31:69:@39748.4]
  wire [15:0] _T_91322; // @[Mux.scala 31:69:@39749.4]
  wire [15:0] _T_91323; // @[Mux.scala 31:69:@39750.4]
  wire [15:0] _T_91324; // @[Mux.scala 31:69:@39751.4]
  wire [15:0] _T_91325; // @[Mux.scala 31:69:@39752.4]
  wire [15:0] _T_91326; // @[Mux.scala 31:69:@39753.4]
  wire [15:0] _T_91327; // @[Mux.scala 31:69:@39754.4]
  wire [15:0] _T_91328; // @[Mux.scala 31:69:@39755.4]
  wire [15:0] _T_91329; // @[Mux.scala 31:69:@39756.4]
  wire [15:0] _T_91330; // @[Mux.scala 31:69:@39757.4]
  wire [15:0] _T_91331; // @[Mux.scala 31:69:@39758.4]
  wire [15:0] _T_91332; // @[Mux.scala 31:69:@39759.4]
  wire [15:0] _T_91333; // @[Mux.scala 31:69:@39760.4]
  wire [15:0] _T_91334; // @[Mux.scala 31:69:@39761.4]
  wire [15:0] _T_91335; // @[Mux.scala 31:69:@39762.4]
  wire  _T_91336; // @[OneHot.scala 66:30:@39763.4]
  wire  _T_91337; // @[OneHot.scala 66:30:@39764.4]
  wire  _T_91338; // @[OneHot.scala 66:30:@39765.4]
  wire  _T_91339; // @[OneHot.scala 66:30:@39766.4]
  wire  _T_91340; // @[OneHot.scala 66:30:@39767.4]
  wire  _T_91341; // @[OneHot.scala 66:30:@39768.4]
  wire  _T_91342; // @[OneHot.scala 66:30:@39769.4]
  wire  _T_91343; // @[OneHot.scala 66:30:@39770.4]
  wire  _T_91344; // @[OneHot.scala 66:30:@39771.4]
  wire  _T_91345; // @[OneHot.scala 66:30:@39772.4]
  wire  _T_91346; // @[OneHot.scala 66:30:@39773.4]
  wire  _T_91347; // @[OneHot.scala 66:30:@39774.4]
  wire  _T_91348; // @[OneHot.scala 66:30:@39775.4]
  wire  _T_91349; // @[OneHot.scala 66:30:@39776.4]
  wire  _T_91350; // @[OneHot.scala 66:30:@39777.4]
  wire  _T_91351; // @[OneHot.scala 66:30:@39778.4]
  wire [15:0] _T_91392; // @[Mux.scala 31:69:@39796.4]
  wire [15:0] _T_91393; // @[Mux.scala 31:69:@39797.4]
  wire [15:0] _T_91394; // @[Mux.scala 31:69:@39798.4]
  wire [15:0] _T_91395; // @[Mux.scala 31:69:@39799.4]
  wire [15:0] _T_91396; // @[Mux.scala 31:69:@39800.4]
  wire [15:0] _T_91397; // @[Mux.scala 31:69:@39801.4]
  wire [15:0] _T_91398; // @[Mux.scala 31:69:@39802.4]
  wire [15:0] _T_91399; // @[Mux.scala 31:69:@39803.4]
  wire [15:0] _T_91400; // @[Mux.scala 31:69:@39804.4]
  wire [15:0] _T_91401; // @[Mux.scala 31:69:@39805.4]
  wire [15:0] _T_91402; // @[Mux.scala 31:69:@39806.4]
  wire [15:0] _T_91403; // @[Mux.scala 31:69:@39807.4]
  wire [15:0] _T_91404; // @[Mux.scala 31:69:@39808.4]
  wire [15:0] _T_91405; // @[Mux.scala 31:69:@39809.4]
  wire [15:0] _T_91406; // @[Mux.scala 31:69:@39810.4]
  wire [15:0] _T_91407; // @[Mux.scala 31:69:@39811.4]
  wire  _T_91408; // @[OneHot.scala 66:30:@39812.4]
  wire  _T_91409; // @[OneHot.scala 66:30:@39813.4]
  wire  _T_91410; // @[OneHot.scala 66:30:@39814.4]
  wire  _T_91411; // @[OneHot.scala 66:30:@39815.4]
  wire  _T_91412; // @[OneHot.scala 66:30:@39816.4]
  wire  _T_91413; // @[OneHot.scala 66:30:@39817.4]
  wire  _T_91414; // @[OneHot.scala 66:30:@39818.4]
  wire  _T_91415; // @[OneHot.scala 66:30:@39819.4]
  wire  _T_91416; // @[OneHot.scala 66:30:@39820.4]
  wire  _T_91417; // @[OneHot.scala 66:30:@39821.4]
  wire  _T_91418; // @[OneHot.scala 66:30:@39822.4]
  wire  _T_91419; // @[OneHot.scala 66:30:@39823.4]
  wire  _T_91420; // @[OneHot.scala 66:30:@39824.4]
  wire  _T_91421; // @[OneHot.scala 66:30:@39825.4]
  wire  _T_91422; // @[OneHot.scala 66:30:@39826.4]
  wire  _T_91423; // @[OneHot.scala 66:30:@39827.4]
  wire [15:0] _T_91464; // @[Mux.scala 31:69:@39845.4]
  wire [15:0] _T_91465; // @[Mux.scala 31:69:@39846.4]
  wire [15:0] _T_91466; // @[Mux.scala 31:69:@39847.4]
  wire [15:0] _T_91467; // @[Mux.scala 31:69:@39848.4]
  wire [15:0] _T_91468; // @[Mux.scala 31:69:@39849.4]
  wire [15:0] _T_91469; // @[Mux.scala 31:69:@39850.4]
  wire [15:0] _T_91470; // @[Mux.scala 31:69:@39851.4]
  wire [15:0] _T_91471; // @[Mux.scala 31:69:@39852.4]
  wire [15:0] _T_91472; // @[Mux.scala 31:69:@39853.4]
  wire [15:0] _T_91473; // @[Mux.scala 31:69:@39854.4]
  wire [15:0] _T_91474; // @[Mux.scala 31:69:@39855.4]
  wire [15:0] _T_91475; // @[Mux.scala 31:69:@39856.4]
  wire [15:0] _T_91476; // @[Mux.scala 31:69:@39857.4]
  wire [15:0] _T_91477; // @[Mux.scala 31:69:@39858.4]
  wire [15:0] _T_91478; // @[Mux.scala 31:69:@39859.4]
  wire [15:0] _T_91479; // @[Mux.scala 31:69:@39860.4]
  wire  _T_91480; // @[OneHot.scala 66:30:@39861.4]
  wire  _T_91481; // @[OneHot.scala 66:30:@39862.4]
  wire  _T_91482; // @[OneHot.scala 66:30:@39863.4]
  wire  _T_91483; // @[OneHot.scala 66:30:@39864.4]
  wire  _T_91484; // @[OneHot.scala 66:30:@39865.4]
  wire  _T_91485; // @[OneHot.scala 66:30:@39866.4]
  wire  _T_91486; // @[OneHot.scala 66:30:@39867.4]
  wire  _T_91487; // @[OneHot.scala 66:30:@39868.4]
  wire  _T_91488; // @[OneHot.scala 66:30:@39869.4]
  wire  _T_91489; // @[OneHot.scala 66:30:@39870.4]
  wire  _T_91490; // @[OneHot.scala 66:30:@39871.4]
  wire  _T_91491; // @[OneHot.scala 66:30:@39872.4]
  wire  _T_91492; // @[OneHot.scala 66:30:@39873.4]
  wire  _T_91493; // @[OneHot.scala 66:30:@39874.4]
  wire  _T_91494; // @[OneHot.scala 66:30:@39875.4]
  wire  _T_91495; // @[OneHot.scala 66:30:@39876.4]
  wire [15:0] _T_91536; // @[Mux.scala 31:69:@39894.4]
  wire [15:0] _T_91537; // @[Mux.scala 31:69:@39895.4]
  wire [15:0] _T_91538; // @[Mux.scala 31:69:@39896.4]
  wire [15:0] _T_91539; // @[Mux.scala 31:69:@39897.4]
  wire [15:0] _T_91540; // @[Mux.scala 31:69:@39898.4]
  wire [15:0] _T_91541; // @[Mux.scala 31:69:@39899.4]
  wire [15:0] _T_91542; // @[Mux.scala 31:69:@39900.4]
  wire [15:0] _T_91543; // @[Mux.scala 31:69:@39901.4]
  wire [15:0] _T_91544; // @[Mux.scala 31:69:@39902.4]
  wire [15:0] _T_91545; // @[Mux.scala 31:69:@39903.4]
  wire [15:0] _T_91546; // @[Mux.scala 31:69:@39904.4]
  wire [15:0] _T_91547; // @[Mux.scala 31:69:@39905.4]
  wire [15:0] _T_91548; // @[Mux.scala 31:69:@39906.4]
  wire [15:0] _T_91549; // @[Mux.scala 31:69:@39907.4]
  wire [15:0] _T_91550; // @[Mux.scala 31:69:@39908.4]
  wire [15:0] _T_91551; // @[Mux.scala 31:69:@39909.4]
  wire  _T_91552; // @[OneHot.scala 66:30:@39910.4]
  wire  _T_91553; // @[OneHot.scala 66:30:@39911.4]
  wire  _T_91554; // @[OneHot.scala 66:30:@39912.4]
  wire  _T_91555; // @[OneHot.scala 66:30:@39913.4]
  wire  _T_91556; // @[OneHot.scala 66:30:@39914.4]
  wire  _T_91557; // @[OneHot.scala 66:30:@39915.4]
  wire  _T_91558; // @[OneHot.scala 66:30:@39916.4]
  wire  _T_91559; // @[OneHot.scala 66:30:@39917.4]
  wire  _T_91560; // @[OneHot.scala 66:30:@39918.4]
  wire  _T_91561; // @[OneHot.scala 66:30:@39919.4]
  wire  _T_91562; // @[OneHot.scala 66:30:@39920.4]
  wire  _T_91563; // @[OneHot.scala 66:30:@39921.4]
  wire  _T_91564; // @[OneHot.scala 66:30:@39922.4]
  wire  _T_91565; // @[OneHot.scala 66:30:@39923.4]
  wire  _T_91566; // @[OneHot.scala 66:30:@39924.4]
  wire  _T_91567; // @[OneHot.scala 66:30:@39925.4]
  wire [7:0] _T_91632; // @[Mux.scala 19:72:@39949.4]
  wire [15:0] _T_91640; // @[Mux.scala 19:72:@39957.4]
  wire [15:0] _T_91642; // @[Mux.scala 19:72:@39958.4]
  wire [7:0] _T_91649; // @[Mux.scala 19:72:@39965.4]
  wire [15:0] _T_91657; // @[Mux.scala 19:72:@39973.4]
  wire [15:0] _T_91659; // @[Mux.scala 19:72:@39974.4]
  wire [7:0] _T_91666; // @[Mux.scala 19:72:@39981.4]
  wire [15:0] _T_91674; // @[Mux.scala 19:72:@39989.4]
  wire [15:0] _T_91676; // @[Mux.scala 19:72:@39990.4]
  wire [7:0] _T_91683; // @[Mux.scala 19:72:@39997.4]
  wire [15:0] _T_91691; // @[Mux.scala 19:72:@40005.4]
  wire [15:0] _T_91693; // @[Mux.scala 19:72:@40006.4]
  wire [7:0] _T_91700; // @[Mux.scala 19:72:@40013.4]
  wire [15:0] _T_91708; // @[Mux.scala 19:72:@40021.4]
  wire [15:0] _T_91710; // @[Mux.scala 19:72:@40022.4]
  wire [7:0] _T_91717; // @[Mux.scala 19:72:@40029.4]
  wire [15:0] _T_91725; // @[Mux.scala 19:72:@40037.4]
  wire [15:0] _T_91727; // @[Mux.scala 19:72:@40038.4]
  wire [7:0] _T_91734; // @[Mux.scala 19:72:@40045.4]
  wire [15:0] _T_91742; // @[Mux.scala 19:72:@40053.4]
  wire [15:0] _T_91744; // @[Mux.scala 19:72:@40054.4]
  wire [7:0] _T_91751; // @[Mux.scala 19:72:@40061.4]
  wire [15:0] _T_91759; // @[Mux.scala 19:72:@40069.4]
  wire [15:0] _T_91761; // @[Mux.scala 19:72:@40070.4]
  wire [7:0] _T_91768; // @[Mux.scala 19:72:@40077.4]
  wire [15:0] _T_91776; // @[Mux.scala 19:72:@40085.4]
  wire [15:0] _T_91778; // @[Mux.scala 19:72:@40086.4]
  wire [7:0] _T_91785; // @[Mux.scala 19:72:@40093.4]
  wire [15:0] _T_91793; // @[Mux.scala 19:72:@40101.4]
  wire [15:0] _T_91795; // @[Mux.scala 19:72:@40102.4]
  wire [7:0] _T_91802; // @[Mux.scala 19:72:@40109.4]
  wire [15:0] _T_91810; // @[Mux.scala 19:72:@40117.4]
  wire [15:0] _T_91812; // @[Mux.scala 19:72:@40118.4]
  wire [7:0] _T_91819; // @[Mux.scala 19:72:@40125.4]
  wire [15:0] _T_91827; // @[Mux.scala 19:72:@40133.4]
  wire [15:0] _T_91829; // @[Mux.scala 19:72:@40134.4]
  wire [7:0] _T_91836; // @[Mux.scala 19:72:@40141.4]
  wire [15:0] _T_91844; // @[Mux.scala 19:72:@40149.4]
  wire [15:0] _T_91846; // @[Mux.scala 19:72:@40150.4]
  wire [7:0] _T_91853; // @[Mux.scala 19:72:@40157.4]
  wire [15:0] _T_91861; // @[Mux.scala 19:72:@40165.4]
  wire [15:0] _T_91863; // @[Mux.scala 19:72:@40166.4]
  wire [7:0] _T_91870; // @[Mux.scala 19:72:@40173.4]
  wire [15:0] _T_91878; // @[Mux.scala 19:72:@40181.4]
  wire [15:0] _T_91880; // @[Mux.scala 19:72:@40182.4]
  wire [7:0] _T_91887; // @[Mux.scala 19:72:@40189.4]
  wire [15:0] _T_91895; // @[Mux.scala 19:72:@40197.4]
  wire [15:0] _T_91897; // @[Mux.scala 19:72:@40198.4]
  wire [15:0] _T_91898; // @[Mux.scala 19:72:@40199.4]
  wire [15:0] _T_91899; // @[Mux.scala 19:72:@40200.4]
  wire [15:0] _T_91900; // @[Mux.scala 19:72:@40201.4]
  wire [15:0] _T_91901; // @[Mux.scala 19:72:@40202.4]
  wire [15:0] _T_91902; // @[Mux.scala 19:72:@40203.4]
  wire [15:0] _T_91903; // @[Mux.scala 19:72:@40204.4]
  wire [15:0] _T_91904; // @[Mux.scala 19:72:@40205.4]
  wire [15:0] _T_91905; // @[Mux.scala 19:72:@40206.4]
  wire [15:0] _T_91906; // @[Mux.scala 19:72:@40207.4]
  wire [15:0] _T_91907; // @[Mux.scala 19:72:@40208.4]
  wire [15:0] _T_91908; // @[Mux.scala 19:72:@40209.4]
  wire [15:0] _T_91909; // @[Mux.scala 19:72:@40210.4]
  wire [15:0] _T_91910; // @[Mux.scala 19:72:@40211.4]
  wire [15:0] _T_91911; // @[Mux.scala 19:72:@40212.4]
  wire [15:0] _T_91912; // @[Mux.scala 19:72:@40213.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@40217.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@40219.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@40221.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@40223.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@40225.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@40227.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@40229.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@40231.4]
  wire  priorityLoadRequest_8; // @[Mux.scala 19:72:@40233.4]
  wire  priorityLoadRequest_9; // @[Mux.scala 19:72:@40235.4]
  wire  priorityLoadRequest_10; // @[Mux.scala 19:72:@40237.4]
  wire  priorityLoadRequest_11; // @[Mux.scala 19:72:@40239.4]
  wire  priorityLoadRequest_12; // @[Mux.scala 19:72:@40241.4]
  wire  priorityLoadRequest_13; // @[Mux.scala 19:72:@40243.4]
  wire  priorityLoadRequest_14; // @[Mux.scala 19:72:@40245.4]
  wire  priorityLoadRequest_15; // @[Mux.scala 19:72:@40247.4]
  wire  _GEN_1920; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1921; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1922; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1923; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1924; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1925; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1926; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1927; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1928; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1929; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1930; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1931; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1932; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1933; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1934; // @[LoadQueue.scala 208:31:@40267.4]
  wire  _GEN_1935; // @[LoadQueue.scala 208:31:@40267.4]
  wire [7:0] _T_92307; // @[LoadQueue.scala 238:58:@40485.8]
  wire [15:0] _T_92315; // @[LoadQueue.scala 238:58:@40493.8]
  wire [7:0] _T_92322; // @[LoadQueue.scala 238:96:@40500.8]
  wire [15:0] _T_92330; // @[LoadQueue.scala 238:96:@40508.8]
  wire  _T_92331; // @[LoadQueue.scala 238:61:@40509.8]
  wire  _T_92332; // @[LoadQueue.scala 237:64:@40510.8]
  wire  _GEN_1969; // @[LoadQueue.scala 230:110:@40442.6]
  wire  bypassRequest_0; // @[LoadQueue.scala 229:71:@40436.4]
  wire  _GEN_1936; // @[LoadQueue.scala 217:34:@40324.6]
  wire  _GEN_1937; // @[LoadQueue.scala 215:23:@40320.4]
  wire [7:0] _T_92391; // @[LoadQueue.scala 238:58:@40567.8]
  wire [15:0] _T_92399; // @[LoadQueue.scala 238:58:@40575.8]
  wire [7:0] _T_92406; // @[LoadQueue.scala 238:96:@40582.8]
  wire [15:0] _T_92414; // @[LoadQueue.scala 238:96:@40590.8]
  wire  _T_92415; // @[LoadQueue.scala 238:61:@40591.8]
  wire  _T_92416; // @[LoadQueue.scala 237:64:@40592.8]
  wire  _GEN_1973; // @[LoadQueue.scala 230:110:@40524.6]
  wire  bypassRequest_1; // @[LoadQueue.scala 229:71:@40518.4]
  wire  _GEN_1938; // @[LoadQueue.scala 217:34:@40331.6]
  wire  _GEN_1939; // @[LoadQueue.scala 215:23:@40327.4]
  wire [7:0] _T_92475; // @[LoadQueue.scala 238:58:@40649.8]
  wire [15:0] _T_92483; // @[LoadQueue.scala 238:58:@40657.8]
  wire [7:0] _T_92490; // @[LoadQueue.scala 238:96:@40664.8]
  wire [15:0] _T_92498; // @[LoadQueue.scala 238:96:@40672.8]
  wire  _T_92499; // @[LoadQueue.scala 238:61:@40673.8]
  wire  _T_92500; // @[LoadQueue.scala 237:64:@40674.8]
  wire  _GEN_1977; // @[LoadQueue.scala 230:110:@40606.6]
  wire  bypassRequest_2; // @[LoadQueue.scala 229:71:@40600.4]
  wire  _GEN_1940; // @[LoadQueue.scala 217:34:@40338.6]
  wire  _GEN_1941; // @[LoadQueue.scala 215:23:@40334.4]
  wire [7:0] _T_92559; // @[LoadQueue.scala 238:58:@40731.8]
  wire [15:0] _T_92567; // @[LoadQueue.scala 238:58:@40739.8]
  wire [7:0] _T_92574; // @[LoadQueue.scala 238:96:@40746.8]
  wire [15:0] _T_92582; // @[LoadQueue.scala 238:96:@40754.8]
  wire  _T_92583; // @[LoadQueue.scala 238:61:@40755.8]
  wire  _T_92584; // @[LoadQueue.scala 237:64:@40756.8]
  wire  _GEN_1981; // @[LoadQueue.scala 230:110:@40688.6]
  wire  bypassRequest_3; // @[LoadQueue.scala 229:71:@40682.4]
  wire  _GEN_1942; // @[LoadQueue.scala 217:34:@40345.6]
  wire  _GEN_1943; // @[LoadQueue.scala 215:23:@40341.4]
  wire [7:0] _T_92643; // @[LoadQueue.scala 238:58:@40813.8]
  wire [15:0] _T_92651; // @[LoadQueue.scala 238:58:@40821.8]
  wire [7:0] _T_92658; // @[LoadQueue.scala 238:96:@40828.8]
  wire [15:0] _T_92666; // @[LoadQueue.scala 238:96:@40836.8]
  wire  _T_92667; // @[LoadQueue.scala 238:61:@40837.8]
  wire  _T_92668; // @[LoadQueue.scala 237:64:@40838.8]
  wire  _GEN_1985; // @[LoadQueue.scala 230:110:@40770.6]
  wire  bypassRequest_4; // @[LoadQueue.scala 229:71:@40764.4]
  wire  _GEN_1944; // @[LoadQueue.scala 217:34:@40352.6]
  wire  _GEN_1945; // @[LoadQueue.scala 215:23:@40348.4]
  wire [7:0] _T_92727; // @[LoadQueue.scala 238:58:@40895.8]
  wire [15:0] _T_92735; // @[LoadQueue.scala 238:58:@40903.8]
  wire [7:0] _T_92742; // @[LoadQueue.scala 238:96:@40910.8]
  wire [15:0] _T_92750; // @[LoadQueue.scala 238:96:@40918.8]
  wire  _T_92751; // @[LoadQueue.scala 238:61:@40919.8]
  wire  _T_92752; // @[LoadQueue.scala 237:64:@40920.8]
  wire  _GEN_1989; // @[LoadQueue.scala 230:110:@40852.6]
  wire  bypassRequest_5; // @[LoadQueue.scala 229:71:@40846.4]
  wire  _GEN_1946; // @[LoadQueue.scala 217:34:@40359.6]
  wire  _GEN_1947; // @[LoadQueue.scala 215:23:@40355.4]
  wire [7:0] _T_92811; // @[LoadQueue.scala 238:58:@40977.8]
  wire [15:0] _T_92819; // @[LoadQueue.scala 238:58:@40985.8]
  wire [7:0] _T_92826; // @[LoadQueue.scala 238:96:@40992.8]
  wire [15:0] _T_92834; // @[LoadQueue.scala 238:96:@41000.8]
  wire  _T_92835; // @[LoadQueue.scala 238:61:@41001.8]
  wire  _T_92836; // @[LoadQueue.scala 237:64:@41002.8]
  wire  _GEN_1993; // @[LoadQueue.scala 230:110:@40934.6]
  wire  bypassRequest_6; // @[LoadQueue.scala 229:71:@40928.4]
  wire  _GEN_1948; // @[LoadQueue.scala 217:34:@40366.6]
  wire  _GEN_1949; // @[LoadQueue.scala 215:23:@40362.4]
  wire [7:0] _T_92895; // @[LoadQueue.scala 238:58:@41059.8]
  wire [15:0] _T_92903; // @[LoadQueue.scala 238:58:@41067.8]
  wire [7:0] _T_92910; // @[LoadQueue.scala 238:96:@41074.8]
  wire [15:0] _T_92918; // @[LoadQueue.scala 238:96:@41082.8]
  wire  _T_92919; // @[LoadQueue.scala 238:61:@41083.8]
  wire  _T_92920; // @[LoadQueue.scala 237:64:@41084.8]
  wire  _GEN_1997; // @[LoadQueue.scala 230:110:@41016.6]
  wire  bypassRequest_7; // @[LoadQueue.scala 229:71:@41010.4]
  wire  _GEN_1950; // @[LoadQueue.scala 217:34:@40373.6]
  wire  _GEN_1951; // @[LoadQueue.scala 215:23:@40369.4]
  wire [7:0] _T_92979; // @[LoadQueue.scala 238:58:@41141.8]
  wire [15:0] _T_92987; // @[LoadQueue.scala 238:58:@41149.8]
  wire [7:0] _T_92994; // @[LoadQueue.scala 238:96:@41156.8]
  wire [15:0] _T_93002; // @[LoadQueue.scala 238:96:@41164.8]
  wire  _T_93003; // @[LoadQueue.scala 238:61:@41165.8]
  wire  _T_93004; // @[LoadQueue.scala 237:64:@41166.8]
  wire  _GEN_2001; // @[LoadQueue.scala 230:110:@41098.6]
  wire  bypassRequest_8; // @[LoadQueue.scala 229:71:@41092.4]
  wire  _GEN_1952; // @[LoadQueue.scala 217:34:@40380.6]
  wire  _GEN_1953; // @[LoadQueue.scala 215:23:@40376.4]
  wire [7:0] _T_93063; // @[LoadQueue.scala 238:58:@41223.8]
  wire [15:0] _T_93071; // @[LoadQueue.scala 238:58:@41231.8]
  wire [7:0] _T_93078; // @[LoadQueue.scala 238:96:@41238.8]
  wire [15:0] _T_93086; // @[LoadQueue.scala 238:96:@41246.8]
  wire  _T_93087; // @[LoadQueue.scala 238:61:@41247.8]
  wire  _T_93088; // @[LoadQueue.scala 237:64:@41248.8]
  wire  _GEN_2005; // @[LoadQueue.scala 230:110:@41180.6]
  wire  bypassRequest_9; // @[LoadQueue.scala 229:71:@41174.4]
  wire  _GEN_1954; // @[LoadQueue.scala 217:34:@40387.6]
  wire  _GEN_1955; // @[LoadQueue.scala 215:23:@40383.4]
  wire [7:0] _T_93147; // @[LoadQueue.scala 238:58:@41305.8]
  wire [15:0] _T_93155; // @[LoadQueue.scala 238:58:@41313.8]
  wire [7:0] _T_93162; // @[LoadQueue.scala 238:96:@41320.8]
  wire [15:0] _T_93170; // @[LoadQueue.scala 238:96:@41328.8]
  wire  _T_93171; // @[LoadQueue.scala 238:61:@41329.8]
  wire  _T_93172; // @[LoadQueue.scala 237:64:@41330.8]
  wire  _GEN_2009; // @[LoadQueue.scala 230:110:@41262.6]
  wire  bypassRequest_10; // @[LoadQueue.scala 229:71:@41256.4]
  wire  _GEN_1956; // @[LoadQueue.scala 217:34:@40394.6]
  wire  _GEN_1957; // @[LoadQueue.scala 215:23:@40390.4]
  wire [7:0] _T_93231; // @[LoadQueue.scala 238:58:@41387.8]
  wire [15:0] _T_93239; // @[LoadQueue.scala 238:58:@41395.8]
  wire [7:0] _T_93246; // @[LoadQueue.scala 238:96:@41402.8]
  wire [15:0] _T_93254; // @[LoadQueue.scala 238:96:@41410.8]
  wire  _T_93255; // @[LoadQueue.scala 238:61:@41411.8]
  wire  _T_93256; // @[LoadQueue.scala 237:64:@41412.8]
  wire  _GEN_2013; // @[LoadQueue.scala 230:110:@41344.6]
  wire  bypassRequest_11; // @[LoadQueue.scala 229:71:@41338.4]
  wire  _GEN_1958; // @[LoadQueue.scala 217:34:@40401.6]
  wire  _GEN_1959; // @[LoadQueue.scala 215:23:@40397.4]
  wire [7:0] _T_93315; // @[LoadQueue.scala 238:58:@41469.8]
  wire [15:0] _T_93323; // @[LoadQueue.scala 238:58:@41477.8]
  wire [7:0] _T_93330; // @[LoadQueue.scala 238:96:@41484.8]
  wire [15:0] _T_93338; // @[LoadQueue.scala 238:96:@41492.8]
  wire  _T_93339; // @[LoadQueue.scala 238:61:@41493.8]
  wire  _T_93340; // @[LoadQueue.scala 237:64:@41494.8]
  wire  _GEN_2017; // @[LoadQueue.scala 230:110:@41426.6]
  wire  bypassRequest_12; // @[LoadQueue.scala 229:71:@41420.4]
  wire  _GEN_1960; // @[LoadQueue.scala 217:34:@40408.6]
  wire  _GEN_1961; // @[LoadQueue.scala 215:23:@40404.4]
  wire [7:0] _T_93399; // @[LoadQueue.scala 238:58:@41551.8]
  wire [15:0] _T_93407; // @[LoadQueue.scala 238:58:@41559.8]
  wire [7:0] _T_93414; // @[LoadQueue.scala 238:96:@41566.8]
  wire [15:0] _T_93422; // @[LoadQueue.scala 238:96:@41574.8]
  wire  _T_93423; // @[LoadQueue.scala 238:61:@41575.8]
  wire  _T_93424; // @[LoadQueue.scala 237:64:@41576.8]
  wire  _GEN_2021; // @[LoadQueue.scala 230:110:@41508.6]
  wire  bypassRequest_13; // @[LoadQueue.scala 229:71:@41502.4]
  wire  _GEN_1962; // @[LoadQueue.scala 217:34:@40415.6]
  wire  _GEN_1963; // @[LoadQueue.scala 215:23:@40411.4]
  wire [7:0] _T_93483; // @[LoadQueue.scala 238:58:@41633.8]
  wire [15:0] _T_93491; // @[LoadQueue.scala 238:58:@41641.8]
  wire [7:0] _T_93498; // @[LoadQueue.scala 238:96:@41648.8]
  wire [15:0] _T_93506; // @[LoadQueue.scala 238:96:@41656.8]
  wire  _T_93507; // @[LoadQueue.scala 238:61:@41657.8]
  wire  _T_93508; // @[LoadQueue.scala 237:64:@41658.8]
  wire  _GEN_2025; // @[LoadQueue.scala 230:110:@41590.6]
  wire  bypassRequest_14; // @[LoadQueue.scala 229:71:@41584.4]
  wire  _GEN_1964; // @[LoadQueue.scala 217:34:@40422.6]
  wire  _GEN_1965; // @[LoadQueue.scala 215:23:@40418.4]
  wire [7:0] _T_93567; // @[LoadQueue.scala 238:58:@41715.8]
  wire [15:0] _T_93575; // @[LoadQueue.scala 238:58:@41723.8]
  wire [7:0] _T_93582; // @[LoadQueue.scala 238:96:@41730.8]
  wire [15:0] _T_93590; // @[LoadQueue.scala 238:96:@41738.8]
  wire  _T_93591; // @[LoadQueue.scala 238:61:@41739.8]
  wire  _T_93592; // @[LoadQueue.scala 237:64:@41740.8]
  wire  _GEN_2029; // @[LoadQueue.scala 230:110:@41672.6]
  wire  bypassRequest_15; // @[LoadQueue.scala 229:71:@41666.4]
  wire  _GEN_1966; // @[LoadQueue.scala 217:34:@40429.6]
  wire  _GEN_1967; // @[LoadQueue.scala 215:23:@40425.4]
  wire  _T_93596; // @[LoadQueue.scala 247:28:@41746.4]
  wire  _T_93597; // @[LoadQueue.scala 247:28:@41747.4]
  wire  _T_93598; // @[LoadQueue.scala 247:28:@41748.4]
  wire  _T_93599; // @[LoadQueue.scala 247:28:@41749.4]
  wire  _T_93600; // @[LoadQueue.scala 247:28:@41750.4]
  wire  _T_93601; // @[LoadQueue.scala 247:28:@41751.4]
  wire  _T_93602; // @[LoadQueue.scala 247:28:@41752.4]
  wire  _T_93603; // @[LoadQueue.scala 247:28:@41753.4]
  wire  _T_93604; // @[LoadQueue.scala 247:28:@41754.4]
  wire  _T_93605; // @[LoadQueue.scala 247:28:@41755.4]
  wire  _T_93606; // @[LoadQueue.scala 247:28:@41756.4]
  wire  _T_93607; // @[LoadQueue.scala 247:28:@41757.4]
  wire  _T_93608; // @[LoadQueue.scala 247:28:@41758.4]
  wire  _T_93609; // @[LoadQueue.scala 247:28:@41759.4]
  wire  _T_93610; // @[LoadQueue.scala 247:28:@41760.4]
  wire [3:0] _T_93627; // @[Mux.scala 31:69:@41762.6]
  wire [3:0] _T_93628; // @[Mux.scala 31:69:@41763.6]
  wire [3:0] _T_93629; // @[Mux.scala 31:69:@41764.6]
  wire [3:0] _T_93630; // @[Mux.scala 31:69:@41765.6]
  wire [3:0] _T_93631; // @[Mux.scala 31:69:@41766.6]
  wire [3:0] _T_93632; // @[Mux.scala 31:69:@41767.6]
  wire [3:0] _T_93633; // @[Mux.scala 31:69:@41768.6]
  wire [3:0] _T_93634; // @[Mux.scala 31:69:@41769.6]
  wire [3:0] _T_93635; // @[Mux.scala 31:69:@41770.6]
  wire [3:0] _T_93636; // @[Mux.scala 31:69:@41771.6]
  wire [3:0] _T_93637; // @[Mux.scala 31:69:@41772.6]
  wire [3:0] _T_93638; // @[Mux.scala 31:69:@41773.6]
  wire [3:0] _T_93639; // @[Mux.scala 31:69:@41774.6]
  wire [3:0] _T_93640; // @[Mux.scala 31:69:@41775.6]
  wire [3:0] _T_93641; // @[Mux.scala 31:69:@41776.6]
  wire [31:0] _GEN_2033; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2034; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2035; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2036; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2037; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2038; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2039; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2040; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2041; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2042; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2043; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2044; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2045; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2046; // @[LoadQueue.scala 248:24:@41777.6]
  wire [31:0] _GEN_2047; // @[LoadQueue.scala 248:24:@41777.6]
  wire  _T_93649; // @[LoadQueue.scala 261:41:@41788.6]
  wire  _GEN_2050; // @[LoadQueue.scala 261:62:@41789.6]
  wire  _GEN_2051; // @[LoadQueue.scala 259:25:@41784.4]
  wire  _T_93652; // @[LoadQueue.scala 261:41:@41796.6]
  wire  _GEN_2052; // @[LoadQueue.scala 261:62:@41797.6]
  wire  _GEN_2053; // @[LoadQueue.scala 259:25:@41792.4]
  wire  _T_93655; // @[LoadQueue.scala 261:41:@41804.6]
  wire  _GEN_2054; // @[LoadQueue.scala 261:62:@41805.6]
  wire  _GEN_2055; // @[LoadQueue.scala 259:25:@41800.4]
  wire  _T_93658; // @[LoadQueue.scala 261:41:@41812.6]
  wire  _GEN_2056; // @[LoadQueue.scala 261:62:@41813.6]
  wire  _GEN_2057; // @[LoadQueue.scala 259:25:@41808.4]
  wire  _T_93661; // @[LoadQueue.scala 261:41:@41820.6]
  wire  _GEN_2058; // @[LoadQueue.scala 261:62:@41821.6]
  wire  _GEN_2059; // @[LoadQueue.scala 259:25:@41816.4]
  wire  _T_93664; // @[LoadQueue.scala 261:41:@41828.6]
  wire  _GEN_2060; // @[LoadQueue.scala 261:62:@41829.6]
  wire  _GEN_2061; // @[LoadQueue.scala 259:25:@41824.4]
  wire  _T_93667; // @[LoadQueue.scala 261:41:@41836.6]
  wire  _GEN_2062; // @[LoadQueue.scala 261:62:@41837.6]
  wire  _GEN_2063; // @[LoadQueue.scala 259:25:@41832.4]
  wire  _T_93670; // @[LoadQueue.scala 261:41:@41844.6]
  wire  _GEN_2064; // @[LoadQueue.scala 261:62:@41845.6]
  wire  _GEN_2065; // @[LoadQueue.scala 259:25:@41840.4]
  wire  _T_93673; // @[LoadQueue.scala 261:41:@41852.6]
  wire  _GEN_2066; // @[LoadQueue.scala 261:62:@41853.6]
  wire  _GEN_2067; // @[LoadQueue.scala 259:25:@41848.4]
  wire  _T_93676; // @[LoadQueue.scala 261:41:@41860.6]
  wire  _GEN_2068; // @[LoadQueue.scala 261:62:@41861.6]
  wire  _GEN_2069; // @[LoadQueue.scala 259:25:@41856.4]
  wire  _T_93679; // @[LoadQueue.scala 261:41:@41868.6]
  wire  _GEN_2070; // @[LoadQueue.scala 261:62:@41869.6]
  wire  _GEN_2071; // @[LoadQueue.scala 259:25:@41864.4]
  wire  _T_93682; // @[LoadQueue.scala 261:41:@41876.6]
  wire  _GEN_2072; // @[LoadQueue.scala 261:62:@41877.6]
  wire  _GEN_2073; // @[LoadQueue.scala 259:25:@41872.4]
  wire  _T_93685; // @[LoadQueue.scala 261:41:@41884.6]
  wire  _GEN_2074; // @[LoadQueue.scala 261:62:@41885.6]
  wire  _GEN_2075; // @[LoadQueue.scala 259:25:@41880.4]
  wire  _T_93688; // @[LoadQueue.scala 261:41:@41892.6]
  wire  _GEN_2076; // @[LoadQueue.scala 261:62:@41893.6]
  wire  _GEN_2077; // @[LoadQueue.scala 259:25:@41888.4]
  wire  _T_93691; // @[LoadQueue.scala 261:41:@41900.6]
  wire  _GEN_2078; // @[LoadQueue.scala 261:62:@41901.6]
  wire  _GEN_2079; // @[LoadQueue.scala 259:25:@41896.4]
  wire  _T_93694; // @[LoadQueue.scala 261:41:@41908.6]
  wire  _GEN_2080; // @[LoadQueue.scala 261:62:@41909.6]
  wire  _GEN_2081; // @[LoadQueue.scala 259:25:@41904.4]
  wire [31:0] _GEN_2082; // @[LoadQueue.scala 269:44:@41916.6]
  wire [31:0] _GEN_2083; // @[LoadQueue.scala 267:32:@41912.4]
  wire [31:0] _GEN_2084; // @[LoadQueue.scala 269:44:@41923.6]
  wire [31:0] _GEN_2085; // @[LoadQueue.scala 267:32:@41919.4]
  wire [31:0] _GEN_2086; // @[LoadQueue.scala 269:44:@41930.6]
  wire [31:0] _GEN_2087; // @[LoadQueue.scala 267:32:@41926.4]
  wire [31:0] _GEN_2088; // @[LoadQueue.scala 269:44:@41937.6]
  wire [31:0] _GEN_2089; // @[LoadQueue.scala 267:32:@41933.4]
  wire [31:0] _GEN_2090; // @[LoadQueue.scala 269:44:@41944.6]
  wire [31:0] _GEN_2091; // @[LoadQueue.scala 267:32:@41940.4]
  wire [31:0] _GEN_2092; // @[LoadQueue.scala 269:44:@41951.6]
  wire [31:0] _GEN_2093; // @[LoadQueue.scala 267:32:@41947.4]
  wire [31:0] _GEN_2094; // @[LoadQueue.scala 269:44:@41958.6]
  wire [31:0] _GEN_2095; // @[LoadQueue.scala 267:32:@41954.4]
  wire [31:0] _GEN_2096; // @[LoadQueue.scala 269:44:@41965.6]
  wire [31:0] _GEN_2097; // @[LoadQueue.scala 267:32:@41961.4]
  wire [31:0] _GEN_2098; // @[LoadQueue.scala 269:44:@41972.6]
  wire [31:0] _GEN_2099; // @[LoadQueue.scala 267:32:@41968.4]
  wire [31:0] _GEN_2100; // @[LoadQueue.scala 269:44:@41979.6]
  wire [31:0] _GEN_2101; // @[LoadQueue.scala 267:32:@41975.4]
  wire [31:0] _GEN_2102; // @[LoadQueue.scala 269:44:@41986.6]
  wire [31:0] _GEN_2103; // @[LoadQueue.scala 267:32:@41982.4]
  wire [31:0] _GEN_2104; // @[LoadQueue.scala 269:44:@41993.6]
  wire [31:0] _GEN_2105; // @[LoadQueue.scala 267:32:@41989.4]
  wire [31:0] _GEN_2106; // @[LoadQueue.scala 269:44:@42000.6]
  wire [31:0] _GEN_2107; // @[LoadQueue.scala 267:32:@41996.4]
  wire [31:0] _GEN_2108; // @[LoadQueue.scala 269:44:@42007.6]
  wire [31:0] _GEN_2109; // @[LoadQueue.scala 267:32:@42003.4]
  wire [31:0] _GEN_2110; // @[LoadQueue.scala 269:44:@42014.6]
  wire [31:0] _GEN_2111; // @[LoadQueue.scala 267:32:@42010.4]
  wire [31:0] _GEN_2112; // @[LoadQueue.scala 269:44:@42021.6]
  wire [31:0] _GEN_2113; // @[LoadQueue.scala 267:32:@42017.4]
  wire  entriesPorts_0_0; // @[LoadQueue.scala 286:69:@42025.4]
  wire  entriesPorts_0_1; // @[LoadQueue.scala 286:69:@42027.4]
  wire  entriesPorts_0_2; // @[LoadQueue.scala 286:69:@42029.4]
  wire  entriesPorts_0_3; // @[LoadQueue.scala 286:69:@42031.4]
  wire  entriesPorts_0_4; // @[LoadQueue.scala 286:69:@42033.4]
  wire  entriesPorts_0_5; // @[LoadQueue.scala 286:69:@42035.4]
  wire  entriesPorts_0_6; // @[LoadQueue.scala 286:69:@42037.4]
  wire  entriesPorts_0_7; // @[LoadQueue.scala 286:69:@42039.4]
  wire  entriesPorts_0_8; // @[LoadQueue.scala 286:69:@42041.4]
  wire  entriesPorts_0_9; // @[LoadQueue.scala 286:69:@42043.4]
  wire  entriesPorts_0_10; // @[LoadQueue.scala 286:69:@42045.4]
  wire  entriesPorts_0_11; // @[LoadQueue.scala 286:69:@42047.4]
  wire  entriesPorts_0_12; // @[LoadQueue.scala 286:69:@42049.4]
  wire  entriesPorts_0_13; // @[LoadQueue.scala 286:69:@42051.4]
  wire  entriesPorts_0_14; // @[LoadQueue.scala 286:69:@42053.4]
  wire  entriesPorts_0_15; // @[LoadQueue.scala 286:69:@42055.4]
  wire  _T_94179; // @[LoadQueue.scala 298:86:@42059.4]
  wire  _T_94180; // @[LoadQueue.scala 298:83:@42060.4]
  wire  _T_94182; // @[LoadQueue.scala 298:86:@42061.4]
  wire  _T_94183; // @[LoadQueue.scala 298:83:@42062.4]
  wire  _T_94185; // @[LoadQueue.scala 298:86:@42063.4]
  wire  _T_94186; // @[LoadQueue.scala 298:83:@42064.4]
  wire  _T_94188; // @[LoadQueue.scala 298:86:@42065.4]
  wire  _T_94189; // @[LoadQueue.scala 298:83:@42066.4]
  wire  _T_94191; // @[LoadQueue.scala 298:86:@42067.4]
  wire  _T_94192; // @[LoadQueue.scala 298:83:@42068.4]
  wire  _T_94194; // @[LoadQueue.scala 298:86:@42069.4]
  wire  _T_94195; // @[LoadQueue.scala 298:83:@42070.4]
  wire  _T_94197; // @[LoadQueue.scala 298:86:@42071.4]
  wire  _T_94198; // @[LoadQueue.scala 298:83:@42072.4]
  wire  _T_94200; // @[LoadQueue.scala 298:86:@42073.4]
  wire  _T_94201; // @[LoadQueue.scala 298:83:@42074.4]
  wire  _T_94203; // @[LoadQueue.scala 298:86:@42075.4]
  wire  _T_94204; // @[LoadQueue.scala 298:83:@42076.4]
  wire  _T_94206; // @[LoadQueue.scala 298:86:@42077.4]
  wire  _T_94207; // @[LoadQueue.scala 298:83:@42078.4]
  wire  _T_94209; // @[LoadQueue.scala 298:86:@42079.4]
  wire  _T_94210; // @[LoadQueue.scala 298:83:@42080.4]
  wire  _T_94212; // @[LoadQueue.scala 298:86:@42081.4]
  wire  _T_94213; // @[LoadQueue.scala 298:83:@42082.4]
  wire  _T_94215; // @[LoadQueue.scala 298:86:@42083.4]
  wire  _T_94216; // @[LoadQueue.scala 298:83:@42084.4]
  wire  _T_94218; // @[LoadQueue.scala 298:86:@42085.4]
  wire  _T_94219; // @[LoadQueue.scala 298:83:@42086.4]
  wire  _T_94221; // @[LoadQueue.scala 298:86:@42087.4]
  wire  _T_94222; // @[LoadQueue.scala 298:83:@42088.4]
  wire  _T_94224; // @[LoadQueue.scala 298:86:@42089.4]
  wire  _T_94225; // @[LoadQueue.scala 298:83:@42090.4]
  wire [15:0] _T_94308; // @[Mux.scala 31:69:@42144.4]
  wire [15:0] _T_94309; // @[Mux.scala 31:69:@42145.4]
  wire [15:0] _T_94310; // @[Mux.scala 31:69:@42146.4]
  wire [15:0] _T_94311; // @[Mux.scala 31:69:@42147.4]
  wire [15:0] _T_94312; // @[Mux.scala 31:69:@42148.4]
  wire [15:0] _T_94313; // @[Mux.scala 31:69:@42149.4]
  wire [15:0] _T_94314; // @[Mux.scala 31:69:@42150.4]
  wire [15:0] _T_94315; // @[Mux.scala 31:69:@42151.4]
  wire [15:0] _T_94316; // @[Mux.scala 31:69:@42152.4]
  wire [15:0] _T_94317; // @[Mux.scala 31:69:@42153.4]
  wire [15:0] _T_94318; // @[Mux.scala 31:69:@42154.4]
  wire [15:0] _T_94319; // @[Mux.scala 31:69:@42155.4]
  wire [15:0] _T_94320; // @[Mux.scala 31:69:@42156.4]
  wire [15:0] _T_94321; // @[Mux.scala 31:69:@42157.4]
  wire [15:0] _T_94322; // @[Mux.scala 31:69:@42158.4]
  wire [15:0] _T_94323; // @[Mux.scala 31:69:@42159.4]
  wire  _T_94324; // @[OneHot.scala 66:30:@42160.4]
  wire  _T_94325; // @[OneHot.scala 66:30:@42161.4]
  wire  _T_94326; // @[OneHot.scala 66:30:@42162.4]
  wire  _T_94327; // @[OneHot.scala 66:30:@42163.4]
  wire  _T_94328; // @[OneHot.scala 66:30:@42164.4]
  wire  _T_94329; // @[OneHot.scala 66:30:@42165.4]
  wire  _T_94330; // @[OneHot.scala 66:30:@42166.4]
  wire  _T_94331; // @[OneHot.scala 66:30:@42167.4]
  wire  _T_94332; // @[OneHot.scala 66:30:@42168.4]
  wire  _T_94333; // @[OneHot.scala 66:30:@42169.4]
  wire  _T_94334; // @[OneHot.scala 66:30:@42170.4]
  wire  _T_94335; // @[OneHot.scala 66:30:@42171.4]
  wire  _T_94336; // @[OneHot.scala 66:30:@42172.4]
  wire  _T_94337; // @[OneHot.scala 66:30:@42173.4]
  wire  _T_94338; // @[OneHot.scala 66:30:@42174.4]
  wire  _T_94339; // @[OneHot.scala 66:30:@42175.4]
  wire [15:0] _T_94380; // @[Mux.scala 31:69:@42193.4]
  wire [15:0] _T_94381; // @[Mux.scala 31:69:@42194.4]
  wire [15:0] _T_94382; // @[Mux.scala 31:69:@42195.4]
  wire [15:0] _T_94383; // @[Mux.scala 31:69:@42196.4]
  wire [15:0] _T_94384; // @[Mux.scala 31:69:@42197.4]
  wire [15:0] _T_94385; // @[Mux.scala 31:69:@42198.4]
  wire [15:0] _T_94386; // @[Mux.scala 31:69:@42199.4]
  wire [15:0] _T_94387; // @[Mux.scala 31:69:@42200.4]
  wire [15:0] _T_94388; // @[Mux.scala 31:69:@42201.4]
  wire [15:0] _T_94389; // @[Mux.scala 31:69:@42202.4]
  wire [15:0] _T_94390; // @[Mux.scala 31:69:@42203.4]
  wire [15:0] _T_94391; // @[Mux.scala 31:69:@42204.4]
  wire [15:0] _T_94392; // @[Mux.scala 31:69:@42205.4]
  wire [15:0] _T_94393; // @[Mux.scala 31:69:@42206.4]
  wire [15:0] _T_94394; // @[Mux.scala 31:69:@42207.4]
  wire [15:0] _T_94395; // @[Mux.scala 31:69:@42208.4]
  wire  _T_94396; // @[OneHot.scala 66:30:@42209.4]
  wire  _T_94397; // @[OneHot.scala 66:30:@42210.4]
  wire  _T_94398; // @[OneHot.scala 66:30:@42211.4]
  wire  _T_94399; // @[OneHot.scala 66:30:@42212.4]
  wire  _T_94400; // @[OneHot.scala 66:30:@42213.4]
  wire  _T_94401; // @[OneHot.scala 66:30:@42214.4]
  wire  _T_94402; // @[OneHot.scala 66:30:@42215.4]
  wire  _T_94403; // @[OneHot.scala 66:30:@42216.4]
  wire  _T_94404; // @[OneHot.scala 66:30:@42217.4]
  wire  _T_94405; // @[OneHot.scala 66:30:@42218.4]
  wire  _T_94406; // @[OneHot.scala 66:30:@42219.4]
  wire  _T_94407; // @[OneHot.scala 66:30:@42220.4]
  wire  _T_94408; // @[OneHot.scala 66:30:@42221.4]
  wire  _T_94409; // @[OneHot.scala 66:30:@42222.4]
  wire  _T_94410; // @[OneHot.scala 66:30:@42223.4]
  wire  _T_94411; // @[OneHot.scala 66:30:@42224.4]
  wire [15:0] _T_94452; // @[Mux.scala 31:69:@42242.4]
  wire [15:0] _T_94453; // @[Mux.scala 31:69:@42243.4]
  wire [15:0] _T_94454; // @[Mux.scala 31:69:@42244.4]
  wire [15:0] _T_94455; // @[Mux.scala 31:69:@42245.4]
  wire [15:0] _T_94456; // @[Mux.scala 31:69:@42246.4]
  wire [15:0] _T_94457; // @[Mux.scala 31:69:@42247.4]
  wire [15:0] _T_94458; // @[Mux.scala 31:69:@42248.4]
  wire [15:0] _T_94459; // @[Mux.scala 31:69:@42249.4]
  wire [15:0] _T_94460; // @[Mux.scala 31:69:@42250.4]
  wire [15:0] _T_94461; // @[Mux.scala 31:69:@42251.4]
  wire [15:0] _T_94462; // @[Mux.scala 31:69:@42252.4]
  wire [15:0] _T_94463; // @[Mux.scala 31:69:@42253.4]
  wire [15:0] _T_94464; // @[Mux.scala 31:69:@42254.4]
  wire [15:0] _T_94465; // @[Mux.scala 31:69:@42255.4]
  wire [15:0] _T_94466; // @[Mux.scala 31:69:@42256.4]
  wire [15:0] _T_94467; // @[Mux.scala 31:69:@42257.4]
  wire  _T_94468; // @[OneHot.scala 66:30:@42258.4]
  wire  _T_94469; // @[OneHot.scala 66:30:@42259.4]
  wire  _T_94470; // @[OneHot.scala 66:30:@42260.4]
  wire  _T_94471; // @[OneHot.scala 66:30:@42261.4]
  wire  _T_94472; // @[OneHot.scala 66:30:@42262.4]
  wire  _T_94473; // @[OneHot.scala 66:30:@42263.4]
  wire  _T_94474; // @[OneHot.scala 66:30:@42264.4]
  wire  _T_94475; // @[OneHot.scala 66:30:@42265.4]
  wire  _T_94476; // @[OneHot.scala 66:30:@42266.4]
  wire  _T_94477; // @[OneHot.scala 66:30:@42267.4]
  wire  _T_94478; // @[OneHot.scala 66:30:@42268.4]
  wire  _T_94479; // @[OneHot.scala 66:30:@42269.4]
  wire  _T_94480; // @[OneHot.scala 66:30:@42270.4]
  wire  _T_94481; // @[OneHot.scala 66:30:@42271.4]
  wire  _T_94482; // @[OneHot.scala 66:30:@42272.4]
  wire  _T_94483; // @[OneHot.scala 66:30:@42273.4]
  wire [15:0] _T_94524; // @[Mux.scala 31:69:@42291.4]
  wire [15:0] _T_94525; // @[Mux.scala 31:69:@42292.4]
  wire [15:0] _T_94526; // @[Mux.scala 31:69:@42293.4]
  wire [15:0] _T_94527; // @[Mux.scala 31:69:@42294.4]
  wire [15:0] _T_94528; // @[Mux.scala 31:69:@42295.4]
  wire [15:0] _T_94529; // @[Mux.scala 31:69:@42296.4]
  wire [15:0] _T_94530; // @[Mux.scala 31:69:@42297.4]
  wire [15:0] _T_94531; // @[Mux.scala 31:69:@42298.4]
  wire [15:0] _T_94532; // @[Mux.scala 31:69:@42299.4]
  wire [15:0] _T_94533; // @[Mux.scala 31:69:@42300.4]
  wire [15:0] _T_94534; // @[Mux.scala 31:69:@42301.4]
  wire [15:0] _T_94535; // @[Mux.scala 31:69:@42302.4]
  wire [15:0] _T_94536; // @[Mux.scala 31:69:@42303.4]
  wire [15:0] _T_94537; // @[Mux.scala 31:69:@42304.4]
  wire [15:0] _T_94538; // @[Mux.scala 31:69:@42305.4]
  wire [15:0] _T_94539; // @[Mux.scala 31:69:@42306.4]
  wire  _T_94540; // @[OneHot.scala 66:30:@42307.4]
  wire  _T_94541; // @[OneHot.scala 66:30:@42308.4]
  wire  _T_94542; // @[OneHot.scala 66:30:@42309.4]
  wire  _T_94543; // @[OneHot.scala 66:30:@42310.4]
  wire  _T_94544; // @[OneHot.scala 66:30:@42311.4]
  wire  _T_94545; // @[OneHot.scala 66:30:@42312.4]
  wire  _T_94546; // @[OneHot.scala 66:30:@42313.4]
  wire  _T_94547; // @[OneHot.scala 66:30:@42314.4]
  wire  _T_94548; // @[OneHot.scala 66:30:@42315.4]
  wire  _T_94549; // @[OneHot.scala 66:30:@42316.4]
  wire  _T_94550; // @[OneHot.scala 66:30:@42317.4]
  wire  _T_94551; // @[OneHot.scala 66:30:@42318.4]
  wire  _T_94552; // @[OneHot.scala 66:30:@42319.4]
  wire  _T_94553; // @[OneHot.scala 66:30:@42320.4]
  wire  _T_94554; // @[OneHot.scala 66:30:@42321.4]
  wire  _T_94555; // @[OneHot.scala 66:30:@42322.4]
  wire [15:0] _T_94596; // @[Mux.scala 31:69:@42340.4]
  wire [15:0] _T_94597; // @[Mux.scala 31:69:@42341.4]
  wire [15:0] _T_94598; // @[Mux.scala 31:69:@42342.4]
  wire [15:0] _T_94599; // @[Mux.scala 31:69:@42343.4]
  wire [15:0] _T_94600; // @[Mux.scala 31:69:@42344.4]
  wire [15:0] _T_94601; // @[Mux.scala 31:69:@42345.4]
  wire [15:0] _T_94602; // @[Mux.scala 31:69:@42346.4]
  wire [15:0] _T_94603; // @[Mux.scala 31:69:@42347.4]
  wire [15:0] _T_94604; // @[Mux.scala 31:69:@42348.4]
  wire [15:0] _T_94605; // @[Mux.scala 31:69:@42349.4]
  wire [15:0] _T_94606; // @[Mux.scala 31:69:@42350.4]
  wire [15:0] _T_94607; // @[Mux.scala 31:69:@42351.4]
  wire [15:0] _T_94608; // @[Mux.scala 31:69:@42352.4]
  wire [15:0] _T_94609; // @[Mux.scala 31:69:@42353.4]
  wire [15:0] _T_94610; // @[Mux.scala 31:69:@42354.4]
  wire [15:0] _T_94611; // @[Mux.scala 31:69:@42355.4]
  wire  _T_94612; // @[OneHot.scala 66:30:@42356.4]
  wire  _T_94613; // @[OneHot.scala 66:30:@42357.4]
  wire  _T_94614; // @[OneHot.scala 66:30:@42358.4]
  wire  _T_94615; // @[OneHot.scala 66:30:@42359.4]
  wire  _T_94616; // @[OneHot.scala 66:30:@42360.4]
  wire  _T_94617; // @[OneHot.scala 66:30:@42361.4]
  wire  _T_94618; // @[OneHot.scala 66:30:@42362.4]
  wire  _T_94619; // @[OneHot.scala 66:30:@42363.4]
  wire  _T_94620; // @[OneHot.scala 66:30:@42364.4]
  wire  _T_94621; // @[OneHot.scala 66:30:@42365.4]
  wire  _T_94622; // @[OneHot.scala 66:30:@42366.4]
  wire  _T_94623; // @[OneHot.scala 66:30:@42367.4]
  wire  _T_94624; // @[OneHot.scala 66:30:@42368.4]
  wire  _T_94625; // @[OneHot.scala 66:30:@42369.4]
  wire  _T_94626; // @[OneHot.scala 66:30:@42370.4]
  wire  _T_94627; // @[OneHot.scala 66:30:@42371.4]
  wire [15:0] _T_94668; // @[Mux.scala 31:69:@42389.4]
  wire [15:0] _T_94669; // @[Mux.scala 31:69:@42390.4]
  wire [15:0] _T_94670; // @[Mux.scala 31:69:@42391.4]
  wire [15:0] _T_94671; // @[Mux.scala 31:69:@42392.4]
  wire [15:0] _T_94672; // @[Mux.scala 31:69:@42393.4]
  wire [15:0] _T_94673; // @[Mux.scala 31:69:@42394.4]
  wire [15:0] _T_94674; // @[Mux.scala 31:69:@42395.4]
  wire [15:0] _T_94675; // @[Mux.scala 31:69:@42396.4]
  wire [15:0] _T_94676; // @[Mux.scala 31:69:@42397.4]
  wire [15:0] _T_94677; // @[Mux.scala 31:69:@42398.4]
  wire [15:0] _T_94678; // @[Mux.scala 31:69:@42399.4]
  wire [15:0] _T_94679; // @[Mux.scala 31:69:@42400.4]
  wire [15:0] _T_94680; // @[Mux.scala 31:69:@42401.4]
  wire [15:0] _T_94681; // @[Mux.scala 31:69:@42402.4]
  wire [15:0] _T_94682; // @[Mux.scala 31:69:@42403.4]
  wire [15:0] _T_94683; // @[Mux.scala 31:69:@42404.4]
  wire  _T_94684; // @[OneHot.scala 66:30:@42405.4]
  wire  _T_94685; // @[OneHot.scala 66:30:@42406.4]
  wire  _T_94686; // @[OneHot.scala 66:30:@42407.4]
  wire  _T_94687; // @[OneHot.scala 66:30:@42408.4]
  wire  _T_94688; // @[OneHot.scala 66:30:@42409.4]
  wire  _T_94689; // @[OneHot.scala 66:30:@42410.4]
  wire  _T_94690; // @[OneHot.scala 66:30:@42411.4]
  wire  _T_94691; // @[OneHot.scala 66:30:@42412.4]
  wire  _T_94692; // @[OneHot.scala 66:30:@42413.4]
  wire  _T_94693; // @[OneHot.scala 66:30:@42414.4]
  wire  _T_94694; // @[OneHot.scala 66:30:@42415.4]
  wire  _T_94695; // @[OneHot.scala 66:30:@42416.4]
  wire  _T_94696; // @[OneHot.scala 66:30:@42417.4]
  wire  _T_94697; // @[OneHot.scala 66:30:@42418.4]
  wire  _T_94698; // @[OneHot.scala 66:30:@42419.4]
  wire  _T_94699; // @[OneHot.scala 66:30:@42420.4]
  wire [15:0] _T_94740; // @[Mux.scala 31:69:@42438.4]
  wire [15:0] _T_94741; // @[Mux.scala 31:69:@42439.4]
  wire [15:0] _T_94742; // @[Mux.scala 31:69:@42440.4]
  wire [15:0] _T_94743; // @[Mux.scala 31:69:@42441.4]
  wire [15:0] _T_94744; // @[Mux.scala 31:69:@42442.4]
  wire [15:0] _T_94745; // @[Mux.scala 31:69:@42443.4]
  wire [15:0] _T_94746; // @[Mux.scala 31:69:@42444.4]
  wire [15:0] _T_94747; // @[Mux.scala 31:69:@42445.4]
  wire [15:0] _T_94748; // @[Mux.scala 31:69:@42446.4]
  wire [15:0] _T_94749; // @[Mux.scala 31:69:@42447.4]
  wire [15:0] _T_94750; // @[Mux.scala 31:69:@42448.4]
  wire [15:0] _T_94751; // @[Mux.scala 31:69:@42449.4]
  wire [15:0] _T_94752; // @[Mux.scala 31:69:@42450.4]
  wire [15:0] _T_94753; // @[Mux.scala 31:69:@42451.4]
  wire [15:0] _T_94754; // @[Mux.scala 31:69:@42452.4]
  wire [15:0] _T_94755; // @[Mux.scala 31:69:@42453.4]
  wire  _T_94756; // @[OneHot.scala 66:30:@42454.4]
  wire  _T_94757; // @[OneHot.scala 66:30:@42455.4]
  wire  _T_94758; // @[OneHot.scala 66:30:@42456.4]
  wire  _T_94759; // @[OneHot.scala 66:30:@42457.4]
  wire  _T_94760; // @[OneHot.scala 66:30:@42458.4]
  wire  _T_94761; // @[OneHot.scala 66:30:@42459.4]
  wire  _T_94762; // @[OneHot.scala 66:30:@42460.4]
  wire  _T_94763; // @[OneHot.scala 66:30:@42461.4]
  wire  _T_94764; // @[OneHot.scala 66:30:@42462.4]
  wire  _T_94765; // @[OneHot.scala 66:30:@42463.4]
  wire  _T_94766; // @[OneHot.scala 66:30:@42464.4]
  wire  _T_94767; // @[OneHot.scala 66:30:@42465.4]
  wire  _T_94768; // @[OneHot.scala 66:30:@42466.4]
  wire  _T_94769; // @[OneHot.scala 66:30:@42467.4]
  wire  _T_94770; // @[OneHot.scala 66:30:@42468.4]
  wire  _T_94771; // @[OneHot.scala 66:30:@42469.4]
  wire [15:0] _T_94812; // @[Mux.scala 31:69:@42487.4]
  wire [15:0] _T_94813; // @[Mux.scala 31:69:@42488.4]
  wire [15:0] _T_94814; // @[Mux.scala 31:69:@42489.4]
  wire [15:0] _T_94815; // @[Mux.scala 31:69:@42490.4]
  wire [15:0] _T_94816; // @[Mux.scala 31:69:@42491.4]
  wire [15:0] _T_94817; // @[Mux.scala 31:69:@42492.4]
  wire [15:0] _T_94818; // @[Mux.scala 31:69:@42493.4]
  wire [15:0] _T_94819; // @[Mux.scala 31:69:@42494.4]
  wire [15:0] _T_94820; // @[Mux.scala 31:69:@42495.4]
  wire [15:0] _T_94821; // @[Mux.scala 31:69:@42496.4]
  wire [15:0] _T_94822; // @[Mux.scala 31:69:@42497.4]
  wire [15:0] _T_94823; // @[Mux.scala 31:69:@42498.4]
  wire [15:0] _T_94824; // @[Mux.scala 31:69:@42499.4]
  wire [15:0] _T_94825; // @[Mux.scala 31:69:@42500.4]
  wire [15:0] _T_94826; // @[Mux.scala 31:69:@42501.4]
  wire [15:0] _T_94827; // @[Mux.scala 31:69:@42502.4]
  wire  _T_94828; // @[OneHot.scala 66:30:@42503.4]
  wire  _T_94829; // @[OneHot.scala 66:30:@42504.4]
  wire  _T_94830; // @[OneHot.scala 66:30:@42505.4]
  wire  _T_94831; // @[OneHot.scala 66:30:@42506.4]
  wire  _T_94832; // @[OneHot.scala 66:30:@42507.4]
  wire  _T_94833; // @[OneHot.scala 66:30:@42508.4]
  wire  _T_94834; // @[OneHot.scala 66:30:@42509.4]
  wire  _T_94835; // @[OneHot.scala 66:30:@42510.4]
  wire  _T_94836; // @[OneHot.scala 66:30:@42511.4]
  wire  _T_94837; // @[OneHot.scala 66:30:@42512.4]
  wire  _T_94838; // @[OneHot.scala 66:30:@42513.4]
  wire  _T_94839; // @[OneHot.scala 66:30:@42514.4]
  wire  _T_94840; // @[OneHot.scala 66:30:@42515.4]
  wire  _T_94841; // @[OneHot.scala 66:30:@42516.4]
  wire  _T_94842; // @[OneHot.scala 66:30:@42517.4]
  wire  _T_94843; // @[OneHot.scala 66:30:@42518.4]
  wire [15:0] _T_94884; // @[Mux.scala 31:69:@42536.4]
  wire [15:0] _T_94885; // @[Mux.scala 31:69:@42537.4]
  wire [15:0] _T_94886; // @[Mux.scala 31:69:@42538.4]
  wire [15:0] _T_94887; // @[Mux.scala 31:69:@42539.4]
  wire [15:0] _T_94888; // @[Mux.scala 31:69:@42540.4]
  wire [15:0] _T_94889; // @[Mux.scala 31:69:@42541.4]
  wire [15:0] _T_94890; // @[Mux.scala 31:69:@42542.4]
  wire [15:0] _T_94891; // @[Mux.scala 31:69:@42543.4]
  wire [15:0] _T_94892; // @[Mux.scala 31:69:@42544.4]
  wire [15:0] _T_94893; // @[Mux.scala 31:69:@42545.4]
  wire [15:0] _T_94894; // @[Mux.scala 31:69:@42546.4]
  wire [15:0] _T_94895; // @[Mux.scala 31:69:@42547.4]
  wire [15:0] _T_94896; // @[Mux.scala 31:69:@42548.4]
  wire [15:0] _T_94897; // @[Mux.scala 31:69:@42549.4]
  wire [15:0] _T_94898; // @[Mux.scala 31:69:@42550.4]
  wire [15:0] _T_94899; // @[Mux.scala 31:69:@42551.4]
  wire  _T_94900; // @[OneHot.scala 66:30:@42552.4]
  wire  _T_94901; // @[OneHot.scala 66:30:@42553.4]
  wire  _T_94902; // @[OneHot.scala 66:30:@42554.4]
  wire  _T_94903; // @[OneHot.scala 66:30:@42555.4]
  wire  _T_94904; // @[OneHot.scala 66:30:@42556.4]
  wire  _T_94905; // @[OneHot.scala 66:30:@42557.4]
  wire  _T_94906; // @[OneHot.scala 66:30:@42558.4]
  wire  _T_94907; // @[OneHot.scala 66:30:@42559.4]
  wire  _T_94908; // @[OneHot.scala 66:30:@42560.4]
  wire  _T_94909; // @[OneHot.scala 66:30:@42561.4]
  wire  _T_94910; // @[OneHot.scala 66:30:@42562.4]
  wire  _T_94911; // @[OneHot.scala 66:30:@42563.4]
  wire  _T_94912; // @[OneHot.scala 66:30:@42564.4]
  wire  _T_94913; // @[OneHot.scala 66:30:@42565.4]
  wire  _T_94914; // @[OneHot.scala 66:30:@42566.4]
  wire  _T_94915; // @[OneHot.scala 66:30:@42567.4]
  wire [15:0] _T_94956; // @[Mux.scala 31:69:@42585.4]
  wire [15:0] _T_94957; // @[Mux.scala 31:69:@42586.4]
  wire [15:0] _T_94958; // @[Mux.scala 31:69:@42587.4]
  wire [15:0] _T_94959; // @[Mux.scala 31:69:@42588.4]
  wire [15:0] _T_94960; // @[Mux.scala 31:69:@42589.4]
  wire [15:0] _T_94961; // @[Mux.scala 31:69:@42590.4]
  wire [15:0] _T_94962; // @[Mux.scala 31:69:@42591.4]
  wire [15:0] _T_94963; // @[Mux.scala 31:69:@42592.4]
  wire [15:0] _T_94964; // @[Mux.scala 31:69:@42593.4]
  wire [15:0] _T_94965; // @[Mux.scala 31:69:@42594.4]
  wire [15:0] _T_94966; // @[Mux.scala 31:69:@42595.4]
  wire [15:0] _T_94967; // @[Mux.scala 31:69:@42596.4]
  wire [15:0] _T_94968; // @[Mux.scala 31:69:@42597.4]
  wire [15:0] _T_94969; // @[Mux.scala 31:69:@42598.4]
  wire [15:0] _T_94970; // @[Mux.scala 31:69:@42599.4]
  wire [15:0] _T_94971; // @[Mux.scala 31:69:@42600.4]
  wire  _T_94972; // @[OneHot.scala 66:30:@42601.4]
  wire  _T_94973; // @[OneHot.scala 66:30:@42602.4]
  wire  _T_94974; // @[OneHot.scala 66:30:@42603.4]
  wire  _T_94975; // @[OneHot.scala 66:30:@42604.4]
  wire  _T_94976; // @[OneHot.scala 66:30:@42605.4]
  wire  _T_94977; // @[OneHot.scala 66:30:@42606.4]
  wire  _T_94978; // @[OneHot.scala 66:30:@42607.4]
  wire  _T_94979; // @[OneHot.scala 66:30:@42608.4]
  wire  _T_94980; // @[OneHot.scala 66:30:@42609.4]
  wire  _T_94981; // @[OneHot.scala 66:30:@42610.4]
  wire  _T_94982; // @[OneHot.scala 66:30:@42611.4]
  wire  _T_94983; // @[OneHot.scala 66:30:@42612.4]
  wire  _T_94984; // @[OneHot.scala 66:30:@42613.4]
  wire  _T_94985; // @[OneHot.scala 66:30:@42614.4]
  wire  _T_94986; // @[OneHot.scala 66:30:@42615.4]
  wire  _T_94987; // @[OneHot.scala 66:30:@42616.4]
  wire [15:0] _T_95028; // @[Mux.scala 31:69:@42634.4]
  wire [15:0] _T_95029; // @[Mux.scala 31:69:@42635.4]
  wire [15:0] _T_95030; // @[Mux.scala 31:69:@42636.4]
  wire [15:0] _T_95031; // @[Mux.scala 31:69:@42637.4]
  wire [15:0] _T_95032; // @[Mux.scala 31:69:@42638.4]
  wire [15:0] _T_95033; // @[Mux.scala 31:69:@42639.4]
  wire [15:0] _T_95034; // @[Mux.scala 31:69:@42640.4]
  wire [15:0] _T_95035; // @[Mux.scala 31:69:@42641.4]
  wire [15:0] _T_95036; // @[Mux.scala 31:69:@42642.4]
  wire [15:0] _T_95037; // @[Mux.scala 31:69:@42643.4]
  wire [15:0] _T_95038; // @[Mux.scala 31:69:@42644.4]
  wire [15:0] _T_95039; // @[Mux.scala 31:69:@42645.4]
  wire [15:0] _T_95040; // @[Mux.scala 31:69:@42646.4]
  wire [15:0] _T_95041; // @[Mux.scala 31:69:@42647.4]
  wire [15:0] _T_95042; // @[Mux.scala 31:69:@42648.4]
  wire [15:0] _T_95043; // @[Mux.scala 31:69:@42649.4]
  wire  _T_95044; // @[OneHot.scala 66:30:@42650.4]
  wire  _T_95045; // @[OneHot.scala 66:30:@42651.4]
  wire  _T_95046; // @[OneHot.scala 66:30:@42652.4]
  wire  _T_95047; // @[OneHot.scala 66:30:@42653.4]
  wire  _T_95048; // @[OneHot.scala 66:30:@42654.4]
  wire  _T_95049; // @[OneHot.scala 66:30:@42655.4]
  wire  _T_95050; // @[OneHot.scala 66:30:@42656.4]
  wire  _T_95051; // @[OneHot.scala 66:30:@42657.4]
  wire  _T_95052; // @[OneHot.scala 66:30:@42658.4]
  wire  _T_95053; // @[OneHot.scala 66:30:@42659.4]
  wire  _T_95054; // @[OneHot.scala 66:30:@42660.4]
  wire  _T_95055; // @[OneHot.scala 66:30:@42661.4]
  wire  _T_95056; // @[OneHot.scala 66:30:@42662.4]
  wire  _T_95057; // @[OneHot.scala 66:30:@42663.4]
  wire  _T_95058; // @[OneHot.scala 66:30:@42664.4]
  wire  _T_95059; // @[OneHot.scala 66:30:@42665.4]
  wire [15:0] _T_95100; // @[Mux.scala 31:69:@42683.4]
  wire [15:0] _T_95101; // @[Mux.scala 31:69:@42684.4]
  wire [15:0] _T_95102; // @[Mux.scala 31:69:@42685.4]
  wire [15:0] _T_95103; // @[Mux.scala 31:69:@42686.4]
  wire [15:0] _T_95104; // @[Mux.scala 31:69:@42687.4]
  wire [15:0] _T_95105; // @[Mux.scala 31:69:@42688.4]
  wire [15:0] _T_95106; // @[Mux.scala 31:69:@42689.4]
  wire [15:0] _T_95107; // @[Mux.scala 31:69:@42690.4]
  wire [15:0] _T_95108; // @[Mux.scala 31:69:@42691.4]
  wire [15:0] _T_95109; // @[Mux.scala 31:69:@42692.4]
  wire [15:0] _T_95110; // @[Mux.scala 31:69:@42693.4]
  wire [15:0] _T_95111; // @[Mux.scala 31:69:@42694.4]
  wire [15:0] _T_95112; // @[Mux.scala 31:69:@42695.4]
  wire [15:0] _T_95113; // @[Mux.scala 31:69:@42696.4]
  wire [15:0] _T_95114; // @[Mux.scala 31:69:@42697.4]
  wire [15:0] _T_95115; // @[Mux.scala 31:69:@42698.4]
  wire  _T_95116; // @[OneHot.scala 66:30:@42699.4]
  wire  _T_95117; // @[OneHot.scala 66:30:@42700.4]
  wire  _T_95118; // @[OneHot.scala 66:30:@42701.4]
  wire  _T_95119; // @[OneHot.scala 66:30:@42702.4]
  wire  _T_95120; // @[OneHot.scala 66:30:@42703.4]
  wire  _T_95121; // @[OneHot.scala 66:30:@42704.4]
  wire  _T_95122; // @[OneHot.scala 66:30:@42705.4]
  wire  _T_95123; // @[OneHot.scala 66:30:@42706.4]
  wire  _T_95124; // @[OneHot.scala 66:30:@42707.4]
  wire  _T_95125; // @[OneHot.scala 66:30:@42708.4]
  wire  _T_95126; // @[OneHot.scala 66:30:@42709.4]
  wire  _T_95127; // @[OneHot.scala 66:30:@42710.4]
  wire  _T_95128; // @[OneHot.scala 66:30:@42711.4]
  wire  _T_95129; // @[OneHot.scala 66:30:@42712.4]
  wire  _T_95130; // @[OneHot.scala 66:30:@42713.4]
  wire  _T_95131; // @[OneHot.scala 66:30:@42714.4]
  wire [15:0] _T_95172; // @[Mux.scala 31:69:@42732.4]
  wire [15:0] _T_95173; // @[Mux.scala 31:69:@42733.4]
  wire [15:0] _T_95174; // @[Mux.scala 31:69:@42734.4]
  wire [15:0] _T_95175; // @[Mux.scala 31:69:@42735.4]
  wire [15:0] _T_95176; // @[Mux.scala 31:69:@42736.4]
  wire [15:0] _T_95177; // @[Mux.scala 31:69:@42737.4]
  wire [15:0] _T_95178; // @[Mux.scala 31:69:@42738.4]
  wire [15:0] _T_95179; // @[Mux.scala 31:69:@42739.4]
  wire [15:0] _T_95180; // @[Mux.scala 31:69:@42740.4]
  wire [15:0] _T_95181; // @[Mux.scala 31:69:@42741.4]
  wire [15:0] _T_95182; // @[Mux.scala 31:69:@42742.4]
  wire [15:0] _T_95183; // @[Mux.scala 31:69:@42743.4]
  wire [15:0] _T_95184; // @[Mux.scala 31:69:@42744.4]
  wire [15:0] _T_95185; // @[Mux.scala 31:69:@42745.4]
  wire [15:0] _T_95186; // @[Mux.scala 31:69:@42746.4]
  wire [15:0] _T_95187; // @[Mux.scala 31:69:@42747.4]
  wire  _T_95188; // @[OneHot.scala 66:30:@42748.4]
  wire  _T_95189; // @[OneHot.scala 66:30:@42749.4]
  wire  _T_95190; // @[OneHot.scala 66:30:@42750.4]
  wire  _T_95191; // @[OneHot.scala 66:30:@42751.4]
  wire  _T_95192; // @[OneHot.scala 66:30:@42752.4]
  wire  _T_95193; // @[OneHot.scala 66:30:@42753.4]
  wire  _T_95194; // @[OneHot.scala 66:30:@42754.4]
  wire  _T_95195; // @[OneHot.scala 66:30:@42755.4]
  wire  _T_95196; // @[OneHot.scala 66:30:@42756.4]
  wire  _T_95197; // @[OneHot.scala 66:30:@42757.4]
  wire  _T_95198; // @[OneHot.scala 66:30:@42758.4]
  wire  _T_95199; // @[OneHot.scala 66:30:@42759.4]
  wire  _T_95200; // @[OneHot.scala 66:30:@42760.4]
  wire  _T_95201; // @[OneHot.scala 66:30:@42761.4]
  wire  _T_95202; // @[OneHot.scala 66:30:@42762.4]
  wire  _T_95203; // @[OneHot.scala 66:30:@42763.4]
  wire [15:0] _T_95244; // @[Mux.scala 31:69:@42781.4]
  wire [15:0] _T_95245; // @[Mux.scala 31:69:@42782.4]
  wire [15:0] _T_95246; // @[Mux.scala 31:69:@42783.4]
  wire [15:0] _T_95247; // @[Mux.scala 31:69:@42784.4]
  wire [15:0] _T_95248; // @[Mux.scala 31:69:@42785.4]
  wire [15:0] _T_95249; // @[Mux.scala 31:69:@42786.4]
  wire [15:0] _T_95250; // @[Mux.scala 31:69:@42787.4]
  wire [15:0] _T_95251; // @[Mux.scala 31:69:@42788.4]
  wire [15:0] _T_95252; // @[Mux.scala 31:69:@42789.4]
  wire [15:0] _T_95253; // @[Mux.scala 31:69:@42790.4]
  wire [15:0] _T_95254; // @[Mux.scala 31:69:@42791.4]
  wire [15:0] _T_95255; // @[Mux.scala 31:69:@42792.4]
  wire [15:0] _T_95256; // @[Mux.scala 31:69:@42793.4]
  wire [15:0] _T_95257; // @[Mux.scala 31:69:@42794.4]
  wire [15:0] _T_95258; // @[Mux.scala 31:69:@42795.4]
  wire [15:0] _T_95259; // @[Mux.scala 31:69:@42796.4]
  wire  _T_95260; // @[OneHot.scala 66:30:@42797.4]
  wire  _T_95261; // @[OneHot.scala 66:30:@42798.4]
  wire  _T_95262; // @[OneHot.scala 66:30:@42799.4]
  wire  _T_95263; // @[OneHot.scala 66:30:@42800.4]
  wire  _T_95264; // @[OneHot.scala 66:30:@42801.4]
  wire  _T_95265; // @[OneHot.scala 66:30:@42802.4]
  wire  _T_95266; // @[OneHot.scala 66:30:@42803.4]
  wire  _T_95267; // @[OneHot.scala 66:30:@42804.4]
  wire  _T_95268; // @[OneHot.scala 66:30:@42805.4]
  wire  _T_95269; // @[OneHot.scala 66:30:@42806.4]
  wire  _T_95270; // @[OneHot.scala 66:30:@42807.4]
  wire  _T_95271; // @[OneHot.scala 66:30:@42808.4]
  wire  _T_95272; // @[OneHot.scala 66:30:@42809.4]
  wire  _T_95273; // @[OneHot.scala 66:30:@42810.4]
  wire  _T_95274; // @[OneHot.scala 66:30:@42811.4]
  wire  _T_95275; // @[OneHot.scala 66:30:@42812.4]
  wire [15:0] _T_95316; // @[Mux.scala 31:69:@42830.4]
  wire [15:0] _T_95317; // @[Mux.scala 31:69:@42831.4]
  wire [15:0] _T_95318; // @[Mux.scala 31:69:@42832.4]
  wire [15:0] _T_95319; // @[Mux.scala 31:69:@42833.4]
  wire [15:0] _T_95320; // @[Mux.scala 31:69:@42834.4]
  wire [15:0] _T_95321; // @[Mux.scala 31:69:@42835.4]
  wire [15:0] _T_95322; // @[Mux.scala 31:69:@42836.4]
  wire [15:0] _T_95323; // @[Mux.scala 31:69:@42837.4]
  wire [15:0] _T_95324; // @[Mux.scala 31:69:@42838.4]
  wire [15:0] _T_95325; // @[Mux.scala 31:69:@42839.4]
  wire [15:0] _T_95326; // @[Mux.scala 31:69:@42840.4]
  wire [15:0] _T_95327; // @[Mux.scala 31:69:@42841.4]
  wire [15:0] _T_95328; // @[Mux.scala 31:69:@42842.4]
  wire [15:0] _T_95329; // @[Mux.scala 31:69:@42843.4]
  wire [15:0] _T_95330; // @[Mux.scala 31:69:@42844.4]
  wire [15:0] _T_95331; // @[Mux.scala 31:69:@42845.4]
  wire  _T_95332; // @[OneHot.scala 66:30:@42846.4]
  wire  _T_95333; // @[OneHot.scala 66:30:@42847.4]
  wire  _T_95334; // @[OneHot.scala 66:30:@42848.4]
  wire  _T_95335; // @[OneHot.scala 66:30:@42849.4]
  wire  _T_95336; // @[OneHot.scala 66:30:@42850.4]
  wire  _T_95337; // @[OneHot.scala 66:30:@42851.4]
  wire  _T_95338; // @[OneHot.scala 66:30:@42852.4]
  wire  _T_95339; // @[OneHot.scala 66:30:@42853.4]
  wire  _T_95340; // @[OneHot.scala 66:30:@42854.4]
  wire  _T_95341; // @[OneHot.scala 66:30:@42855.4]
  wire  _T_95342; // @[OneHot.scala 66:30:@42856.4]
  wire  _T_95343; // @[OneHot.scala 66:30:@42857.4]
  wire  _T_95344; // @[OneHot.scala 66:30:@42858.4]
  wire  _T_95345; // @[OneHot.scala 66:30:@42859.4]
  wire  _T_95346; // @[OneHot.scala 66:30:@42860.4]
  wire  _T_95347; // @[OneHot.scala 66:30:@42861.4]
  wire [15:0] _T_95388; // @[Mux.scala 31:69:@42879.4]
  wire [15:0] _T_95389; // @[Mux.scala 31:69:@42880.4]
  wire [15:0] _T_95390; // @[Mux.scala 31:69:@42881.4]
  wire [15:0] _T_95391; // @[Mux.scala 31:69:@42882.4]
  wire [15:0] _T_95392; // @[Mux.scala 31:69:@42883.4]
  wire [15:0] _T_95393; // @[Mux.scala 31:69:@42884.4]
  wire [15:0] _T_95394; // @[Mux.scala 31:69:@42885.4]
  wire [15:0] _T_95395; // @[Mux.scala 31:69:@42886.4]
  wire [15:0] _T_95396; // @[Mux.scala 31:69:@42887.4]
  wire [15:0] _T_95397; // @[Mux.scala 31:69:@42888.4]
  wire [15:0] _T_95398; // @[Mux.scala 31:69:@42889.4]
  wire [15:0] _T_95399; // @[Mux.scala 31:69:@42890.4]
  wire [15:0] _T_95400; // @[Mux.scala 31:69:@42891.4]
  wire [15:0] _T_95401; // @[Mux.scala 31:69:@42892.4]
  wire [15:0] _T_95402; // @[Mux.scala 31:69:@42893.4]
  wire [15:0] _T_95403; // @[Mux.scala 31:69:@42894.4]
  wire  _T_95404; // @[OneHot.scala 66:30:@42895.4]
  wire  _T_95405; // @[OneHot.scala 66:30:@42896.4]
  wire  _T_95406; // @[OneHot.scala 66:30:@42897.4]
  wire  _T_95407; // @[OneHot.scala 66:30:@42898.4]
  wire  _T_95408; // @[OneHot.scala 66:30:@42899.4]
  wire  _T_95409; // @[OneHot.scala 66:30:@42900.4]
  wire  _T_95410; // @[OneHot.scala 66:30:@42901.4]
  wire  _T_95411; // @[OneHot.scala 66:30:@42902.4]
  wire  _T_95412; // @[OneHot.scala 66:30:@42903.4]
  wire  _T_95413; // @[OneHot.scala 66:30:@42904.4]
  wire  _T_95414; // @[OneHot.scala 66:30:@42905.4]
  wire  _T_95415; // @[OneHot.scala 66:30:@42906.4]
  wire  _T_95416; // @[OneHot.scala 66:30:@42907.4]
  wire  _T_95417; // @[OneHot.scala 66:30:@42908.4]
  wire  _T_95418; // @[OneHot.scala 66:30:@42909.4]
  wire  _T_95419; // @[OneHot.scala 66:30:@42910.4]
  wire [7:0] _T_95484; // @[Mux.scala 19:72:@42934.4]
  wire [15:0] _T_95492; // @[Mux.scala 19:72:@42942.4]
  wire [15:0] _T_95494; // @[Mux.scala 19:72:@42943.4]
  wire [7:0] _T_95501; // @[Mux.scala 19:72:@42950.4]
  wire [15:0] _T_95509; // @[Mux.scala 19:72:@42958.4]
  wire [15:0] _T_95511; // @[Mux.scala 19:72:@42959.4]
  wire [7:0] _T_95518; // @[Mux.scala 19:72:@42966.4]
  wire [15:0] _T_95526; // @[Mux.scala 19:72:@42974.4]
  wire [15:0] _T_95528; // @[Mux.scala 19:72:@42975.4]
  wire [7:0] _T_95535; // @[Mux.scala 19:72:@42982.4]
  wire [15:0] _T_95543; // @[Mux.scala 19:72:@42990.4]
  wire [15:0] _T_95545; // @[Mux.scala 19:72:@42991.4]
  wire [7:0] _T_95552; // @[Mux.scala 19:72:@42998.4]
  wire [15:0] _T_95560; // @[Mux.scala 19:72:@43006.4]
  wire [15:0] _T_95562; // @[Mux.scala 19:72:@43007.4]
  wire [7:0] _T_95569; // @[Mux.scala 19:72:@43014.4]
  wire [15:0] _T_95577; // @[Mux.scala 19:72:@43022.4]
  wire [15:0] _T_95579; // @[Mux.scala 19:72:@43023.4]
  wire [7:0] _T_95586; // @[Mux.scala 19:72:@43030.4]
  wire [15:0] _T_95594; // @[Mux.scala 19:72:@43038.4]
  wire [15:0] _T_95596; // @[Mux.scala 19:72:@43039.4]
  wire [7:0] _T_95603; // @[Mux.scala 19:72:@43046.4]
  wire [15:0] _T_95611; // @[Mux.scala 19:72:@43054.4]
  wire [15:0] _T_95613; // @[Mux.scala 19:72:@43055.4]
  wire [7:0] _T_95620; // @[Mux.scala 19:72:@43062.4]
  wire [15:0] _T_95628; // @[Mux.scala 19:72:@43070.4]
  wire [15:0] _T_95630; // @[Mux.scala 19:72:@43071.4]
  wire [7:0] _T_95637; // @[Mux.scala 19:72:@43078.4]
  wire [15:0] _T_95645; // @[Mux.scala 19:72:@43086.4]
  wire [15:0] _T_95647; // @[Mux.scala 19:72:@43087.4]
  wire [7:0] _T_95654; // @[Mux.scala 19:72:@43094.4]
  wire [15:0] _T_95662; // @[Mux.scala 19:72:@43102.4]
  wire [15:0] _T_95664; // @[Mux.scala 19:72:@43103.4]
  wire [7:0] _T_95671; // @[Mux.scala 19:72:@43110.4]
  wire [15:0] _T_95679; // @[Mux.scala 19:72:@43118.4]
  wire [15:0] _T_95681; // @[Mux.scala 19:72:@43119.4]
  wire [7:0] _T_95688; // @[Mux.scala 19:72:@43126.4]
  wire [15:0] _T_95696; // @[Mux.scala 19:72:@43134.4]
  wire [15:0] _T_95698; // @[Mux.scala 19:72:@43135.4]
  wire [7:0] _T_95705; // @[Mux.scala 19:72:@43142.4]
  wire [15:0] _T_95713; // @[Mux.scala 19:72:@43150.4]
  wire [15:0] _T_95715; // @[Mux.scala 19:72:@43151.4]
  wire [7:0] _T_95722; // @[Mux.scala 19:72:@43158.4]
  wire [15:0] _T_95730; // @[Mux.scala 19:72:@43166.4]
  wire [15:0] _T_95732; // @[Mux.scala 19:72:@43167.4]
  wire [7:0] _T_95739; // @[Mux.scala 19:72:@43174.4]
  wire [15:0] _T_95747; // @[Mux.scala 19:72:@43182.4]
  wire [15:0] _T_95749; // @[Mux.scala 19:72:@43183.4]
  wire [15:0] _T_95750; // @[Mux.scala 19:72:@43184.4]
  wire [15:0] _T_95751; // @[Mux.scala 19:72:@43185.4]
  wire [15:0] _T_95752; // @[Mux.scala 19:72:@43186.4]
  wire [15:0] _T_95753; // @[Mux.scala 19:72:@43187.4]
  wire [15:0] _T_95754; // @[Mux.scala 19:72:@43188.4]
  wire [15:0] _T_95755; // @[Mux.scala 19:72:@43189.4]
  wire [15:0] _T_95756; // @[Mux.scala 19:72:@43190.4]
  wire [15:0] _T_95757; // @[Mux.scala 19:72:@43191.4]
  wire [15:0] _T_95758; // @[Mux.scala 19:72:@43192.4]
  wire [15:0] _T_95759; // @[Mux.scala 19:72:@43193.4]
  wire [15:0] _T_95760; // @[Mux.scala 19:72:@43194.4]
  wire [15:0] _T_95761; // @[Mux.scala 19:72:@43195.4]
  wire [15:0] _T_95762; // @[Mux.scala 19:72:@43196.4]
  wire [15:0] _T_95763; // @[Mux.scala 19:72:@43197.4]
  wire [15:0] _T_95764; // @[Mux.scala 19:72:@43198.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@43202.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@43204.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@43206.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@43208.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@43210.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@43212.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@43214.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@43216.4]
  wire  inputPriorityPorts_0_8; // @[Mux.scala 19:72:@43218.4]
  wire  inputPriorityPorts_0_9; // @[Mux.scala 19:72:@43220.4]
  wire  inputPriorityPorts_0_10; // @[Mux.scala 19:72:@43222.4]
  wire  inputPriorityPorts_0_11; // @[Mux.scala 19:72:@43224.4]
  wire  inputPriorityPorts_0_12; // @[Mux.scala 19:72:@43226.4]
  wire  inputPriorityPorts_0_13; // @[Mux.scala 19:72:@43228.4]
  wire  inputPriorityPorts_0_14; // @[Mux.scala 19:72:@43230.4]
  wire  inputPriorityPorts_0_15; // @[Mux.scala 19:72:@43232.4]
  wire [15:0] _T_95966; // @[Mux.scala 31:69:@43286.4]
  wire [15:0] _T_95967; // @[Mux.scala 31:69:@43287.4]
  wire [15:0] _T_95968; // @[Mux.scala 31:69:@43288.4]
  wire [15:0] _T_95969; // @[Mux.scala 31:69:@43289.4]
  wire [15:0] _T_95970; // @[Mux.scala 31:69:@43290.4]
  wire [15:0] _T_95971; // @[Mux.scala 31:69:@43291.4]
  wire [15:0] _T_95972; // @[Mux.scala 31:69:@43292.4]
  wire [15:0] _T_95973; // @[Mux.scala 31:69:@43293.4]
  wire [15:0] _T_95974; // @[Mux.scala 31:69:@43294.4]
  wire [15:0] _T_95975; // @[Mux.scala 31:69:@43295.4]
  wire [15:0] _T_95976; // @[Mux.scala 31:69:@43296.4]
  wire [15:0] _T_95977; // @[Mux.scala 31:69:@43297.4]
  wire [15:0] _T_95978; // @[Mux.scala 31:69:@43298.4]
  wire [15:0] _T_95979; // @[Mux.scala 31:69:@43299.4]
  wire [15:0] _T_95980; // @[Mux.scala 31:69:@43300.4]
  wire [15:0] _T_95981; // @[Mux.scala 31:69:@43301.4]
  wire  _T_95982; // @[OneHot.scala 66:30:@43302.4]
  wire  _T_95983; // @[OneHot.scala 66:30:@43303.4]
  wire  _T_95984; // @[OneHot.scala 66:30:@43304.4]
  wire  _T_95985; // @[OneHot.scala 66:30:@43305.4]
  wire  _T_95986; // @[OneHot.scala 66:30:@43306.4]
  wire  _T_95987; // @[OneHot.scala 66:30:@43307.4]
  wire  _T_95988; // @[OneHot.scala 66:30:@43308.4]
  wire  _T_95989; // @[OneHot.scala 66:30:@43309.4]
  wire  _T_95990; // @[OneHot.scala 66:30:@43310.4]
  wire  _T_95991; // @[OneHot.scala 66:30:@43311.4]
  wire  _T_95992; // @[OneHot.scala 66:30:@43312.4]
  wire  _T_95993; // @[OneHot.scala 66:30:@43313.4]
  wire  _T_95994; // @[OneHot.scala 66:30:@43314.4]
  wire  _T_95995; // @[OneHot.scala 66:30:@43315.4]
  wire  _T_95996; // @[OneHot.scala 66:30:@43316.4]
  wire  _T_95997; // @[OneHot.scala 66:30:@43317.4]
  wire [15:0] _T_96038; // @[Mux.scala 31:69:@43335.4]
  wire [15:0] _T_96039; // @[Mux.scala 31:69:@43336.4]
  wire [15:0] _T_96040; // @[Mux.scala 31:69:@43337.4]
  wire [15:0] _T_96041; // @[Mux.scala 31:69:@43338.4]
  wire [15:0] _T_96042; // @[Mux.scala 31:69:@43339.4]
  wire [15:0] _T_96043; // @[Mux.scala 31:69:@43340.4]
  wire [15:0] _T_96044; // @[Mux.scala 31:69:@43341.4]
  wire [15:0] _T_96045; // @[Mux.scala 31:69:@43342.4]
  wire [15:0] _T_96046; // @[Mux.scala 31:69:@43343.4]
  wire [15:0] _T_96047; // @[Mux.scala 31:69:@43344.4]
  wire [15:0] _T_96048; // @[Mux.scala 31:69:@43345.4]
  wire [15:0] _T_96049; // @[Mux.scala 31:69:@43346.4]
  wire [15:0] _T_96050; // @[Mux.scala 31:69:@43347.4]
  wire [15:0] _T_96051; // @[Mux.scala 31:69:@43348.4]
  wire [15:0] _T_96052; // @[Mux.scala 31:69:@43349.4]
  wire [15:0] _T_96053; // @[Mux.scala 31:69:@43350.4]
  wire  _T_96054; // @[OneHot.scala 66:30:@43351.4]
  wire  _T_96055; // @[OneHot.scala 66:30:@43352.4]
  wire  _T_96056; // @[OneHot.scala 66:30:@43353.4]
  wire  _T_96057; // @[OneHot.scala 66:30:@43354.4]
  wire  _T_96058; // @[OneHot.scala 66:30:@43355.4]
  wire  _T_96059; // @[OneHot.scala 66:30:@43356.4]
  wire  _T_96060; // @[OneHot.scala 66:30:@43357.4]
  wire  _T_96061; // @[OneHot.scala 66:30:@43358.4]
  wire  _T_96062; // @[OneHot.scala 66:30:@43359.4]
  wire  _T_96063; // @[OneHot.scala 66:30:@43360.4]
  wire  _T_96064; // @[OneHot.scala 66:30:@43361.4]
  wire  _T_96065; // @[OneHot.scala 66:30:@43362.4]
  wire  _T_96066; // @[OneHot.scala 66:30:@43363.4]
  wire  _T_96067; // @[OneHot.scala 66:30:@43364.4]
  wire  _T_96068; // @[OneHot.scala 66:30:@43365.4]
  wire  _T_96069; // @[OneHot.scala 66:30:@43366.4]
  wire [15:0] _T_96110; // @[Mux.scala 31:69:@43384.4]
  wire [15:0] _T_96111; // @[Mux.scala 31:69:@43385.4]
  wire [15:0] _T_96112; // @[Mux.scala 31:69:@43386.4]
  wire [15:0] _T_96113; // @[Mux.scala 31:69:@43387.4]
  wire [15:0] _T_96114; // @[Mux.scala 31:69:@43388.4]
  wire [15:0] _T_96115; // @[Mux.scala 31:69:@43389.4]
  wire [15:0] _T_96116; // @[Mux.scala 31:69:@43390.4]
  wire [15:0] _T_96117; // @[Mux.scala 31:69:@43391.4]
  wire [15:0] _T_96118; // @[Mux.scala 31:69:@43392.4]
  wire [15:0] _T_96119; // @[Mux.scala 31:69:@43393.4]
  wire [15:0] _T_96120; // @[Mux.scala 31:69:@43394.4]
  wire [15:0] _T_96121; // @[Mux.scala 31:69:@43395.4]
  wire [15:0] _T_96122; // @[Mux.scala 31:69:@43396.4]
  wire [15:0] _T_96123; // @[Mux.scala 31:69:@43397.4]
  wire [15:0] _T_96124; // @[Mux.scala 31:69:@43398.4]
  wire [15:0] _T_96125; // @[Mux.scala 31:69:@43399.4]
  wire  _T_96126; // @[OneHot.scala 66:30:@43400.4]
  wire  _T_96127; // @[OneHot.scala 66:30:@43401.4]
  wire  _T_96128; // @[OneHot.scala 66:30:@43402.4]
  wire  _T_96129; // @[OneHot.scala 66:30:@43403.4]
  wire  _T_96130; // @[OneHot.scala 66:30:@43404.4]
  wire  _T_96131; // @[OneHot.scala 66:30:@43405.4]
  wire  _T_96132; // @[OneHot.scala 66:30:@43406.4]
  wire  _T_96133; // @[OneHot.scala 66:30:@43407.4]
  wire  _T_96134; // @[OneHot.scala 66:30:@43408.4]
  wire  _T_96135; // @[OneHot.scala 66:30:@43409.4]
  wire  _T_96136; // @[OneHot.scala 66:30:@43410.4]
  wire  _T_96137; // @[OneHot.scala 66:30:@43411.4]
  wire  _T_96138; // @[OneHot.scala 66:30:@43412.4]
  wire  _T_96139; // @[OneHot.scala 66:30:@43413.4]
  wire  _T_96140; // @[OneHot.scala 66:30:@43414.4]
  wire  _T_96141; // @[OneHot.scala 66:30:@43415.4]
  wire [15:0] _T_96182; // @[Mux.scala 31:69:@43433.4]
  wire [15:0] _T_96183; // @[Mux.scala 31:69:@43434.4]
  wire [15:0] _T_96184; // @[Mux.scala 31:69:@43435.4]
  wire [15:0] _T_96185; // @[Mux.scala 31:69:@43436.4]
  wire [15:0] _T_96186; // @[Mux.scala 31:69:@43437.4]
  wire [15:0] _T_96187; // @[Mux.scala 31:69:@43438.4]
  wire [15:0] _T_96188; // @[Mux.scala 31:69:@43439.4]
  wire [15:0] _T_96189; // @[Mux.scala 31:69:@43440.4]
  wire [15:0] _T_96190; // @[Mux.scala 31:69:@43441.4]
  wire [15:0] _T_96191; // @[Mux.scala 31:69:@43442.4]
  wire [15:0] _T_96192; // @[Mux.scala 31:69:@43443.4]
  wire [15:0] _T_96193; // @[Mux.scala 31:69:@43444.4]
  wire [15:0] _T_96194; // @[Mux.scala 31:69:@43445.4]
  wire [15:0] _T_96195; // @[Mux.scala 31:69:@43446.4]
  wire [15:0] _T_96196; // @[Mux.scala 31:69:@43447.4]
  wire [15:0] _T_96197; // @[Mux.scala 31:69:@43448.4]
  wire  _T_96198; // @[OneHot.scala 66:30:@43449.4]
  wire  _T_96199; // @[OneHot.scala 66:30:@43450.4]
  wire  _T_96200; // @[OneHot.scala 66:30:@43451.4]
  wire  _T_96201; // @[OneHot.scala 66:30:@43452.4]
  wire  _T_96202; // @[OneHot.scala 66:30:@43453.4]
  wire  _T_96203; // @[OneHot.scala 66:30:@43454.4]
  wire  _T_96204; // @[OneHot.scala 66:30:@43455.4]
  wire  _T_96205; // @[OneHot.scala 66:30:@43456.4]
  wire  _T_96206; // @[OneHot.scala 66:30:@43457.4]
  wire  _T_96207; // @[OneHot.scala 66:30:@43458.4]
  wire  _T_96208; // @[OneHot.scala 66:30:@43459.4]
  wire  _T_96209; // @[OneHot.scala 66:30:@43460.4]
  wire  _T_96210; // @[OneHot.scala 66:30:@43461.4]
  wire  _T_96211; // @[OneHot.scala 66:30:@43462.4]
  wire  _T_96212; // @[OneHot.scala 66:30:@43463.4]
  wire  _T_96213; // @[OneHot.scala 66:30:@43464.4]
  wire [15:0] _T_96254; // @[Mux.scala 31:69:@43482.4]
  wire [15:0] _T_96255; // @[Mux.scala 31:69:@43483.4]
  wire [15:0] _T_96256; // @[Mux.scala 31:69:@43484.4]
  wire [15:0] _T_96257; // @[Mux.scala 31:69:@43485.4]
  wire [15:0] _T_96258; // @[Mux.scala 31:69:@43486.4]
  wire [15:0] _T_96259; // @[Mux.scala 31:69:@43487.4]
  wire [15:0] _T_96260; // @[Mux.scala 31:69:@43488.4]
  wire [15:0] _T_96261; // @[Mux.scala 31:69:@43489.4]
  wire [15:0] _T_96262; // @[Mux.scala 31:69:@43490.4]
  wire [15:0] _T_96263; // @[Mux.scala 31:69:@43491.4]
  wire [15:0] _T_96264; // @[Mux.scala 31:69:@43492.4]
  wire [15:0] _T_96265; // @[Mux.scala 31:69:@43493.4]
  wire [15:0] _T_96266; // @[Mux.scala 31:69:@43494.4]
  wire [15:0] _T_96267; // @[Mux.scala 31:69:@43495.4]
  wire [15:0] _T_96268; // @[Mux.scala 31:69:@43496.4]
  wire [15:0] _T_96269; // @[Mux.scala 31:69:@43497.4]
  wire  _T_96270; // @[OneHot.scala 66:30:@43498.4]
  wire  _T_96271; // @[OneHot.scala 66:30:@43499.4]
  wire  _T_96272; // @[OneHot.scala 66:30:@43500.4]
  wire  _T_96273; // @[OneHot.scala 66:30:@43501.4]
  wire  _T_96274; // @[OneHot.scala 66:30:@43502.4]
  wire  _T_96275; // @[OneHot.scala 66:30:@43503.4]
  wire  _T_96276; // @[OneHot.scala 66:30:@43504.4]
  wire  _T_96277; // @[OneHot.scala 66:30:@43505.4]
  wire  _T_96278; // @[OneHot.scala 66:30:@43506.4]
  wire  _T_96279; // @[OneHot.scala 66:30:@43507.4]
  wire  _T_96280; // @[OneHot.scala 66:30:@43508.4]
  wire  _T_96281; // @[OneHot.scala 66:30:@43509.4]
  wire  _T_96282; // @[OneHot.scala 66:30:@43510.4]
  wire  _T_96283; // @[OneHot.scala 66:30:@43511.4]
  wire  _T_96284; // @[OneHot.scala 66:30:@43512.4]
  wire  _T_96285; // @[OneHot.scala 66:30:@43513.4]
  wire [15:0] _T_96326; // @[Mux.scala 31:69:@43531.4]
  wire [15:0] _T_96327; // @[Mux.scala 31:69:@43532.4]
  wire [15:0] _T_96328; // @[Mux.scala 31:69:@43533.4]
  wire [15:0] _T_96329; // @[Mux.scala 31:69:@43534.4]
  wire [15:0] _T_96330; // @[Mux.scala 31:69:@43535.4]
  wire [15:0] _T_96331; // @[Mux.scala 31:69:@43536.4]
  wire [15:0] _T_96332; // @[Mux.scala 31:69:@43537.4]
  wire [15:0] _T_96333; // @[Mux.scala 31:69:@43538.4]
  wire [15:0] _T_96334; // @[Mux.scala 31:69:@43539.4]
  wire [15:0] _T_96335; // @[Mux.scala 31:69:@43540.4]
  wire [15:0] _T_96336; // @[Mux.scala 31:69:@43541.4]
  wire [15:0] _T_96337; // @[Mux.scala 31:69:@43542.4]
  wire [15:0] _T_96338; // @[Mux.scala 31:69:@43543.4]
  wire [15:0] _T_96339; // @[Mux.scala 31:69:@43544.4]
  wire [15:0] _T_96340; // @[Mux.scala 31:69:@43545.4]
  wire [15:0] _T_96341; // @[Mux.scala 31:69:@43546.4]
  wire  _T_96342; // @[OneHot.scala 66:30:@43547.4]
  wire  _T_96343; // @[OneHot.scala 66:30:@43548.4]
  wire  _T_96344; // @[OneHot.scala 66:30:@43549.4]
  wire  _T_96345; // @[OneHot.scala 66:30:@43550.4]
  wire  _T_96346; // @[OneHot.scala 66:30:@43551.4]
  wire  _T_96347; // @[OneHot.scala 66:30:@43552.4]
  wire  _T_96348; // @[OneHot.scala 66:30:@43553.4]
  wire  _T_96349; // @[OneHot.scala 66:30:@43554.4]
  wire  _T_96350; // @[OneHot.scala 66:30:@43555.4]
  wire  _T_96351; // @[OneHot.scala 66:30:@43556.4]
  wire  _T_96352; // @[OneHot.scala 66:30:@43557.4]
  wire  _T_96353; // @[OneHot.scala 66:30:@43558.4]
  wire  _T_96354; // @[OneHot.scala 66:30:@43559.4]
  wire  _T_96355; // @[OneHot.scala 66:30:@43560.4]
  wire  _T_96356; // @[OneHot.scala 66:30:@43561.4]
  wire  _T_96357; // @[OneHot.scala 66:30:@43562.4]
  wire [15:0] _T_96398; // @[Mux.scala 31:69:@43580.4]
  wire [15:0] _T_96399; // @[Mux.scala 31:69:@43581.4]
  wire [15:0] _T_96400; // @[Mux.scala 31:69:@43582.4]
  wire [15:0] _T_96401; // @[Mux.scala 31:69:@43583.4]
  wire [15:0] _T_96402; // @[Mux.scala 31:69:@43584.4]
  wire [15:0] _T_96403; // @[Mux.scala 31:69:@43585.4]
  wire [15:0] _T_96404; // @[Mux.scala 31:69:@43586.4]
  wire [15:0] _T_96405; // @[Mux.scala 31:69:@43587.4]
  wire [15:0] _T_96406; // @[Mux.scala 31:69:@43588.4]
  wire [15:0] _T_96407; // @[Mux.scala 31:69:@43589.4]
  wire [15:0] _T_96408; // @[Mux.scala 31:69:@43590.4]
  wire [15:0] _T_96409; // @[Mux.scala 31:69:@43591.4]
  wire [15:0] _T_96410; // @[Mux.scala 31:69:@43592.4]
  wire [15:0] _T_96411; // @[Mux.scala 31:69:@43593.4]
  wire [15:0] _T_96412; // @[Mux.scala 31:69:@43594.4]
  wire [15:0] _T_96413; // @[Mux.scala 31:69:@43595.4]
  wire  _T_96414; // @[OneHot.scala 66:30:@43596.4]
  wire  _T_96415; // @[OneHot.scala 66:30:@43597.4]
  wire  _T_96416; // @[OneHot.scala 66:30:@43598.4]
  wire  _T_96417; // @[OneHot.scala 66:30:@43599.4]
  wire  _T_96418; // @[OneHot.scala 66:30:@43600.4]
  wire  _T_96419; // @[OneHot.scala 66:30:@43601.4]
  wire  _T_96420; // @[OneHot.scala 66:30:@43602.4]
  wire  _T_96421; // @[OneHot.scala 66:30:@43603.4]
  wire  _T_96422; // @[OneHot.scala 66:30:@43604.4]
  wire  _T_96423; // @[OneHot.scala 66:30:@43605.4]
  wire  _T_96424; // @[OneHot.scala 66:30:@43606.4]
  wire  _T_96425; // @[OneHot.scala 66:30:@43607.4]
  wire  _T_96426; // @[OneHot.scala 66:30:@43608.4]
  wire  _T_96427; // @[OneHot.scala 66:30:@43609.4]
  wire  _T_96428; // @[OneHot.scala 66:30:@43610.4]
  wire  _T_96429; // @[OneHot.scala 66:30:@43611.4]
  wire [15:0] _T_96470; // @[Mux.scala 31:69:@43629.4]
  wire [15:0] _T_96471; // @[Mux.scala 31:69:@43630.4]
  wire [15:0] _T_96472; // @[Mux.scala 31:69:@43631.4]
  wire [15:0] _T_96473; // @[Mux.scala 31:69:@43632.4]
  wire [15:0] _T_96474; // @[Mux.scala 31:69:@43633.4]
  wire [15:0] _T_96475; // @[Mux.scala 31:69:@43634.4]
  wire [15:0] _T_96476; // @[Mux.scala 31:69:@43635.4]
  wire [15:0] _T_96477; // @[Mux.scala 31:69:@43636.4]
  wire [15:0] _T_96478; // @[Mux.scala 31:69:@43637.4]
  wire [15:0] _T_96479; // @[Mux.scala 31:69:@43638.4]
  wire [15:0] _T_96480; // @[Mux.scala 31:69:@43639.4]
  wire [15:0] _T_96481; // @[Mux.scala 31:69:@43640.4]
  wire [15:0] _T_96482; // @[Mux.scala 31:69:@43641.4]
  wire [15:0] _T_96483; // @[Mux.scala 31:69:@43642.4]
  wire [15:0] _T_96484; // @[Mux.scala 31:69:@43643.4]
  wire [15:0] _T_96485; // @[Mux.scala 31:69:@43644.4]
  wire  _T_96486; // @[OneHot.scala 66:30:@43645.4]
  wire  _T_96487; // @[OneHot.scala 66:30:@43646.4]
  wire  _T_96488; // @[OneHot.scala 66:30:@43647.4]
  wire  _T_96489; // @[OneHot.scala 66:30:@43648.4]
  wire  _T_96490; // @[OneHot.scala 66:30:@43649.4]
  wire  _T_96491; // @[OneHot.scala 66:30:@43650.4]
  wire  _T_96492; // @[OneHot.scala 66:30:@43651.4]
  wire  _T_96493; // @[OneHot.scala 66:30:@43652.4]
  wire  _T_96494; // @[OneHot.scala 66:30:@43653.4]
  wire  _T_96495; // @[OneHot.scala 66:30:@43654.4]
  wire  _T_96496; // @[OneHot.scala 66:30:@43655.4]
  wire  _T_96497; // @[OneHot.scala 66:30:@43656.4]
  wire  _T_96498; // @[OneHot.scala 66:30:@43657.4]
  wire  _T_96499; // @[OneHot.scala 66:30:@43658.4]
  wire  _T_96500; // @[OneHot.scala 66:30:@43659.4]
  wire  _T_96501; // @[OneHot.scala 66:30:@43660.4]
  wire [15:0] _T_96542; // @[Mux.scala 31:69:@43678.4]
  wire [15:0] _T_96543; // @[Mux.scala 31:69:@43679.4]
  wire [15:0] _T_96544; // @[Mux.scala 31:69:@43680.4]
  wire [15:0] _T_96545; // @[Mux.scala 31:69:@43681.4]
  wire [15:0] _T_96546; // @[Mux.scala 31:69:@43682.4]
  wire [15:0] _T_96547; // @[Mux.scala 31:69:@43683.4]
  wire [15:0] _T_96548; // @[Mux.scala 31:69:@43684.4]
  wire [15:0] _T_96549; // @[Mux.scala 31:69:@43685.4]
  wire [15:0] _T_96550; // @[Mux.scala 31:69:@43686.4]
  wire [15:0] _T_96551; // @[Mux.scala 31:69:@43687.4]
  wire [15:0] _T_96552; // @[Mux.scala 31:69:@43688.4]
  wire [15:0] _T_96553; // @[Mux.scala 31:69:@43689.4]
  wire [15:0] _T_96554; // @[Mux.scala 31:69:@43690.4]
  wire [15:0] _T_96555; // @[Mux.scala 31:69:@43691.4]
  wire [15:0] _T_96556; // @[Mux.scala 31:69:@43692.4]
  wire [15:0] _T_96557; // @[Mux.scala 31:69:@43693.4]
  wire  _T_96558; // @[OneHot.scala 66:30:@43694.4]
  wire  _T_96559; // @[OneHot.scala 66:30:@43695.4]
  wire  _T_96560; // @[OneHot.scala 66:30:@43696.4]
  wire  _T_96561; // @[OneHot.scala 66:30:@43697.4]
  wire  _T_96562; // @[OneHot.scala 66:30:@43698.4]
  wire  _T_96563; // @[OneHot.scala 66:30:@43699.4]
  wire  _T_96564; // @[OneHot.scala 66:30:@43700.4]
  wire  _T_96565; // @[OneHot.scala 66:30:@43701.4]
  wire  _T_96566; // @[OneHot.scala 66:30:@43702.4]
  wire  _T_96567; // @[OneHot.scala 66:30:@43703.4]
  wire  _T_96568; // @[OneHot.scala 66:30:@43704.4]
  wire  _T_96569; // @[OneHot.scala 66:30:@43705.4]
  wire  _T_96570; // @[OneHot.scala 66:30:@43706.4]
  wire  _T_96571; // @[OneHot.scala 66:30:@43707.4]
  wire  _T_96572; // @[OneHot.scala 66:30:@43708.4]
  wire  _T_96573; // @[OneHot.scala 66:30:@43709.4]
  wire [15:0] _T_96614; // @[Mux.scala 31:69:@43727.4]
  wire [15:0] _T_96615; // @[Mux.scala 31:69:@43728.4]
  wire [15:0] _T_96616; // @[Mux.scala 31:69:@43729.4]
  wire [15:0] _T_96617; // @[Mux.scala 31:69:@43730.4]
  wire [15:0] _T_96618; // @[Mux.scala 31:69:@43731.4]
  wire [15:0] _T_96619; // @[Mux.scala 31:69:@43732.4]
  wire [15:0] _T_96620; // @[Mux.scala 31:69:@43733.4]
  wire [15:0] _T_96621; // @[Mux.scala 31:69:@43734.4]
  wire [15:0] _T_96622; // @[Mux.scala 31:69:@43735.4]
  wire [15:0] _T_96623; // @[Mux.scala 31:69:@43736.4]
  wire [15:0] _T_96624; // @[Mux.scala 31:69:@43737.4]
  wire [15:0] _T_96625; // @[Mux.scala 31:69:@43738.4]
  wire [15:0] _T_96626; // @[Mux.scala 31:69:@43739.4]
  wire [15:0] _T_96627; // @[Mux.scala 31:69:@43740.4]
  wire [15:0] _T_96628; // @[Mux.scala 31:69:@43741.4]
  wire [15:0] _T_96629; // @[Mux.scala 31:69:@43742.4]
  wire  _T_96630; // @[OneHot.scala 66:30:@43743.4]
  wire  _T_96631; // @[OneHot.scala 66:30:@43744.4]
  wire  _T_96632; // @[OneHot.scala 66:30:@43745.4]
  wire  _T_96633; // @[OneHot.scala 66:30:@43746.4]
  wire  _T_96634; // @[OneHot.scala 66:30:@43747.4]
  wire  _T_96635; // @[OneHot.scala 66:30:@43748.4]
  wire  _T_96636; // @[OneHot.scala 66:30:@43749.4]
  wire  _T_96637; // @[OneHot.scala 66:30:@43750.4]
  wire  _T_96638; // @[OneHot.scala 66:30:@43751.4]
  wire  _T_96639; // @[OneHot.scala 66:30:@43752.4]
  wire  _T_96640; // @[OneHot.scala 66:30:@43753.4]
  wire  _T_96641; // @[OneHot.scala 66:30:@43754.4]
  wire  _T_96642; // @[OneHot.scala 66:30:@43755.4]
  wire  _T_96643; // @[OneHot.scala 66:30:@43756.4]
  wire  _T_96644; // @[OneHot.scala 66:30:@43757.4]
  wire  _T_96645; // @[OneHot.scala 66:30:@43758.4]
  wire [15:0] _T_96686; // @[Mux.scala 31:69:@43776.4]
  wire [15:0] _T_96687; // @[Mux.scala 31:69:@43777.4]
  wire [15:0] _T_96688; // @[Mux.scala 31:69:@43778.4]
  wire [15:0] _T_96689; // @[Mux.scala 31:69:@43779.4]
  wire [15:0] _T_96690; // @[Mux.scala 31:69:@43780.4]
  wire [15:0] _T_96691; // @[Mux.scala 31:69:@43781.4]
  wire [15:0] _T_96692; // @[Mux.scala 31:69:@43782.4]
  wire [15:0] _T_96693; // @[Mux.scala 31:69:@43783.4]
  wire [15:0] _T_96694; // @[Mux.scala 31:69:@43784.4]
  wire [15:0] _T_96695; // @[Mux.scala 31:69:@43785.4]
  wire [15:0] _T_96696; // @[Mux.scala 31:69:@43786.4]
  wire [15:0] _T_96697; // @[Mux.scala 31:69:@43787.4]
  wire [15:0] _T_96698; // @[Mux.scala 31:69:@43788.4]
  wire [15:0] _T_96699; // @[Mux.scala 31:69:@43789.4]
  wire [15:0] _T_96700; // @[Mux.scala 31:69:@43790.4]
  wire [15:0] _T_96701; // @[Mux.scala 31:69:@43791.4]
  wire  _T_96702; // @[OneHot.scala 66:30:@43792.4]
  wire  _T_96703; // @[OneHot.scala 66:30:@43793.4]
  wire  _T_96704; // @[OneHot.scala 66:30:@43794.4]
  wire  _T_96705; // @[OneHot.scala 66:30:@43795.4]
  wire  _T_96706; // @[OneHot.scala 66:30:@43796.4]
  wire  _T_96707; // @[OneHot.scala 66:30:@43797.4]
  wire  _T_96708; // @[OneHot.scala 66:30:@43798.4]
  wire  _T_96709; // @[OneHot.scala 66:30:@43799.4]
  wire  _T_96710; // @[OneHot.scala 66:30:@43800.4]
  wire  _T_96711; // @[OneHot.scala 66:30:@43801.4]
  wire  _T_96712; // @[OneHot.scala 66:30:@43802.4]
  wire  _T_96713; // @[OneHot.scala 66:30:@43803.4]
  wire  _T_96714; // @[OneHot.scala 66:30:@43804.4]
  wire  _T_96715; // @[OneHot.scala 66:30:@43805.4]
  wire  _T_96716; // @[OneHot.scala 66:30:@43806.4]
  wire  _T_96717; // @[OneHot.scala 66:30:@43807.4]
  wire [15:0] _T_96758; // @[Mux.scala 31:69:@43825.4]
  wire [15:0] _T_96759; // @[Mux.scala 31:69:@43826.4]
  wire [15:0] _T_96760; // @[Mux.scala 31:69:@43827.4]
  wire [15:0] _T_96761; // @[Mux.scala 31:69:@43828.4]
  wire [15:0] _T_96762; // @[Mux.scala 31:69:@43829.4]
  wire [15:0] _T_96763; // @[Mux.scala 31:69:@43830.4]
  wire [15:0] _T_96764; // @[Mux.scala 31:69:@43831.4]
  wire [15:0] _T_96765; // @[Mux.scala 31:69:@43832.4]
  wire [15:0] _T_96766; // @[Mux.scala 31:69:@43833.4]
  wire [15:0] _T_96767; // @[Mux.scala 31:69:@43834.4]
  wire [15:0] _T_96768; // @[Mux.scala 31:69:@43835.4]
  wire [15:0] _T_96769; // @[Mux.scala 31:69:@43836.4]
  wire [15:0] _T_96770; // @[Mux.scala 31:69:@43837.4]
  wire [15:0] _T_96771; // @[Mux.scala 31:69:@43838.4]
  wire [15:0] _T_96772; // @[Mux.scala 31:69:@43839.4]
  wire [15:0] _T_96773; // @[Mux.scala 31:69:@43840.4]
  wire  _T_96774; // @[OneHot.scala 66:30:@43841.4]
  wire  _T_96775; // @[OneHot.scala 66:30:@43842.4]
  wire  _T_96776; // @[OneHot.scala 66:30:@43843.4]
  wire  _T_96777; // @[OneHot.scala 66:30:@43844.4]
  wire  _T_96778; // @[OneHot.scala 66:30:@43845.4]
  wire  _T_96779; // @[OneHot.scala 66:30:@43846.4]
  wire  _T_96780; // @[OneHot.scala 66:30:@43847.4]
  wire  _T_96781; // @[OneHot.scala 66:30:@43848.4]
  wire  _T_96782; // @[OneHot.scala 66:30:@43849.4]
  wire  _T_96783; // @[OneHot.scala 66:30:@43850.4]
  wire  _T_96784; // @[OneHot.scala 66:30:@43851.4]
  wire  _T_96785; // @[OneHot.scala 66:30:@43852.4]
  wire  _T_96786; // @[OneHot.scala 66:30:@43853.4]
  wire  _T_96787; // @[OneHot.scala 66:30:@43854.4]
  wire  _T_96788; // @[OneHot.scala 66:30:@43855.4]
  wire  _T_96789; // @[OneHot.scala 66:30:@43856.4]
  wire [15:0] _T_96830; // @[Mux.scala 31:69:@43874.4]
  wire [15:0] _T_96831; // @[Mux.scala 31:69:@43875.4]
  wire [15:0] _T_96832; // @[Mux.scala 31:69:@43876.4]
  wire [15:0] _T_96833; // @[Mux.scala 31:69:@43877.4]
  wire [15:0] _T_96834; // @[Mux.scala 31:69:@43878.4]
  wire [15:0] _T_96835; // @[Mux.scala 31:69:@43879.4]
  wire [15:0] _T_96836; // @[Mux.scala 31:69:@43880.4]
  wire [15:0] _T_96837; // @[Mux.scala 31:69:@43881.4]
  wire [15:0] _T_96838; // @[Mux.scala 31:69:@43882.4]
  wire [15:0] _T_96839; // @[Mux.scala 31:69:@43883.4]
  wire [15:0] _T_96840; // @[Mux.scala 31:69:@43884.4]
  wire [15:0] _T_96841; // @[Mux.scala 31:69:@43885.4]
  wire [15:0] _T_96842; // @[Mux.scala 31:69:@43886.4]
  wire [15:0] _T_96843; // @[Mux.scala 31:69:@43887.4]
  wire [15:0] _T_96844; // @[Mux.scala 31:69:@43888.4]
  wire [15:0] _T_96845; // @[Mux.scala 31:69:@43889.4]
  wire  _T_96846; // @[OneHot.scala 66:30:@43890.4]
  wire  _T_96847; // @[OneHot.scala 66:30:@43891.4]
  wire  _T_96848; // @[OneHot.scala 66:30:@43892.4]
  wire  _T_96849; // @[OneHot.scala 66:30:@43893.4]
  wire  _T_96850; // @[OneHot.scala 66:30:@43894.4]
  wire  _T_96851; // @[OneHot.scala 66:30:@43895.4]
  wire  _T_96852; // @[OneHot.scala 66:30:@43896.4]
  wire  _T_96853; // @[OneHot.scala 66:30:@43897.4]
  wire  _T_96854; // @[OneHot.scala 66:30:@43898.4]
  wire  _T_96855; // @[OneHot.scala 66:30:@43899.4]
  wire  _T_96856; // @[OneHot.scala 66:30:@43900.4]
  wire  _T_96857; // @[OneHot.scala 66:30:@43901.4]
  wire  _T_96858; // @[OneHot.scala 66:30:@43902.4]
  wire  _T_96859; // @[OneHot.scala 66:30:@43903.4]
  wire  _T_96860; // @[OneHot.scala 66:30:@43904.4]
  wire  _T_96861; // @[OneHot.scala 66:30:@43905.4]
  wire [15:0] _T_96902; // @[Mux.scala 31:69:@43923.4]
  wire [15:0] _T_96903; // @[Mux.scala 31:69:@43924.4]
  wire [15:0] _T_96904; // @[Mux.scala 31:69:@43925.4]
  wire [15:0] _T_96905; // @[Mux.scala 31:69:@43926.4]
  wire [15:0] _T_96906; // @[Mux.scala 31:69:@43927.4]
  wire [15:0] _T_96907; // @[Mux.scala 31:69:@43928.4]
  wire [15:0] _T_96908; // @[Mux.scala 31:69:@43929.4]
  wire [15:0] _T_96909; // @[Mux.scala 31:69:@43930.4]
  wire [15:0] _T_96910; // @[Mux.scala 31:69:@43931.4]
  wire [15:0] _T_96911; // @[Mux.scala 31:69:@43932.4]
  wire [15:0] _T_96912; // @[Mux.scala 31:69:@43933.4]
  wire [15:0] _T_96913; // @[Mux.scala 31:69:@43934.4]
  wire [15:0] _T_96914; // @[Mux.scala 31:69:@43935.4]
  wire [15:0] _T_96915; // @[Mux.scala 31:69:@43936.4]
  wire [15:0] _T_96916; // @[Mux.scala 31:69:@43937.4]
  wire [15:0] _T_96917; // @[Mux.scala 31:69:@43938.4]
  wire  _T_96918; // @[OneHot.scala 66:30:@43939.4]
  wire  _T_96919; // @[OneHot.scala 66:30:@43940.4]
  wire  _T_96920; // @[OneHot.scala 66:30:@43941.4]
  wire  _T_96921; // @[OneHot.scala 66:30:@43942.4]
  wire  _T_96922; // @[OneHot.scala 66:30:@43943.4]
  wire  _T_96923; // @[OneHot.scala 66:30:@43944.4]
  wire  _T_96924; // @[OneHot.scala 66:30:@43945.4]
  wire  _T_96925; // @[OneHot.scala 66:30:@43946.4]
  wire  _T_96926; // @[OneHot.scala 66:30:@43947.4]
  wire  _T_96927; // @[OneHot.scala 66:30:@43948.4]
  wire  _T_96928; // @[OneHot.scala 66:30:@43949.4]
  wire  _T_96929; // @[OneHot.scala 66:30:@43950.4]
  wire  _T_96930; // @[OneHot.scala 66:30:@43951.4]
  wire  _T_96931; // @[OneHot.scala 66:30:@43952.4]
  wire  _T_96932; // @[OneHot.scala 66:30:@43953.4]
  wire  _T_96933; // @[OneHot.scala 66:30:@43954.4]
  wire [15:0] _T_96974; // @[Mux.scala 31:69:@43972.4]
  wire [15:0] _T_96975; // @[Mux.scala 31:69:@43973.4]
  wire [15:0] _T_96976; // @[Mux.scala 31:69:@43974.4]
  wire [15:0] _T_96977; // @[Mux.scala 31:69:@43975.4]
  wire [15:0] _T_96978; // @[Mux.scala 31:69:@43976.4]
  wire [15:0] _T_96979; // @[Mux.scala 31:69:@43977.4]
  wire [15:0] _T_96980; // @[Mux.scala 31:69:@43978.4]
  wire [15:0] _T_96981; // @[Mux.scala 31:69:@43979.4]
  wire [15:0] _T_96982; // @[Mux.scala 31:69:@43980.4]
  wire [15:0] _T_96983; // @[Mux.scala 31:69:@43981.4]
  wire [15:0] _T_96984; // @[Mux.scala 31:69:@43982.4]
  wire [15:0] _T_96985; // @[Mux.scala 31:69:@43983.4]
  wire [15:0] _T_96986; // @[Mux.scala 31:69:@43984.4]
  wire [15:0] _T_96987; // @[Mux.scala 31:69:@43985.4]
  wire [15:0] _T_96988; // @[Mux.scala 31:69:@43986.4]
  wire [15:0] _T_96989; // @[Mux.scala 31:69:@43987.4]
  wire  _T_96990; // @[OneHot.scala 66:30:@43988.4]
  wire  _T_96991; // @[OneHot.scala 66:30:@43989.4]
  wire  _T_96992; // @[OneHot.scala 66:30:@43990.4]
  wire  _T_96993; // @[OneHot.scala 66:30:@43991.4]
  wire  _T_96994; // @[OneHot.scala 66:30:@43992.4]
  wire  _T_96995; // @[OneHot.scala 66:30:@43993.4]
  wire  _T_96996; // @[OneHot.scala 66:30:@43994.4]
  wire  _T_96997; // @[OneHot.scala 66:30:@43995.4]
  wire  _T_96998; // @[OneHot.scala 66:30:@43996.4]
  wire  _T_96999; // @[OneHot.scala 66:30:@43997.4]
  wire  _T_97000; // @[OneHot.scala 66:30:@43998.4]
  wire  _T_97001; // @[OneHot.scala 66:30:@43999.4]
  wire  _T_97002; // @[OneHot.scala 66:30:@44000.4]
  wire  _T_97003; // @[OneHot.scala 66:30:@44001.4]
  wire  _T_97004; // @[OneHot.scala 66:30:@44002.4]
  wire  _T_97005; // @[OneHot.scala 66:30:@44003.4]
  wire [15:0] _T_97046; // @[Mux.scala 31:69:@44021.4]
  wire [15:0] _T_97047; // @[Mux.scala 31:69:@44022.4]
  wire [15:0] _T_97048; // @[Mux.scala 31:69:@44023.4]
  wire [15:0] _T_97049; // @[Mux.scala 31:69:@44024.4]
  wire [15:0] _T_97050; // @[Mux.scala 31:69:@44025.4]
  wire [15:0] _T_97051; // @[Mux.scala 31:69:@44026.4]
  wire [15:0] _T_97052; // @[Mux.scala 31:69:@44027.4]
  wire [15:0] _T_97053; // @[Mux.scala 31:69:@44028.4]
  wire [15:0] _T_97054; // @[Mux.scala 31:69:@44029.4]
  wire [15:0] _T_97055; // @[Mux.scala 31:69:@44030.4]
  wire [15:0] _T_97056; // @[Mux.scala 31:69:@44031.4]
  wire [15:0] _T_97057; // @[Mux.scala 31:69:@44032.4]
  wire [15:0] _T_97058; // @[Mux.scala 31:69:@44033.4]
  wire [15:0] _T_97059; // @[Mux.scala 31:69:@44034.4]
  wire [15:0] _T_97060; // @[Mux.scala 31:69:@44035.4]
  wire [15:0] _T_97061; // @[Mux.scala 31:69:@44036.4]
  wire  _T_97062; // @[OneHot.scala 66:30:@44037.4]
  wire  _T_97063; // @[OneHot.scala 66:30:@44038.4]
  wire  _T_97064; // @[OneHot.scala 66:30:@44039.4]
  wire  _T_97065; // @[OneHot.scala 66:30:@44040.4]
  wire  _T_97066; // @[OneHot.scala 66:30:@44041.4]
  wire  _T_97067; // @[OneHot.scala 66:30:@44042.4]
  wire  _T_97068; // @[OneHot.scala 66:30:@44043.4]
  wire  _T_97069; // @[OneHot.scala 66:30:@44044.4]
  wire  _T_97070; // @[OneHot.scala 66:30:@44045.4]
  wire  _T_97071; // @[OneHot.scala 66:30:@44046.4]
  wire  _T_97072; // @[OneHot.scala 66:30:@44047.4]
  wire  _T_97073; // @[OneHot.scala 66:30:@44048.4]
  wire  _T_97074; // @[OneHot.scala 66:30:@44049.4]
  wire  _T_97075; // @[OneHot.scala 66:30:@44050.4]
  wire  _T_97076; // @[OneHot.scala 66:30:@44051.4]
  wire  _T_97077; // @[OneHot.scala 66:30:@44052.4]
  wire [7:0] _T_97142; // @[Mux.scala 19:72:@44076.4]
  wire [15:0] _T_97150; // @[Mux.scala 19:72:@44084.4]
  wire [15:0] _T_97152; // @[Mux.scala 19:72:@44085.4]
  wire [7:0] _T_97159; // @[Mux.scala 19:72:@44092.4]
  wire [15:0] _T_97167; // @[Mux.scala 19:72:@44100.4]
  wire [15:0] _T_97169; // @[Mux.scala 19:72:@44101.4]
  wire [7:0] _T_97176; // @[Mux.scala 19:72:@44108.4]
  wire [15:0] _T_97184; // @[Mux.scala 19:72:@44116.4]
  wire [15:0] _T_97186; // @[Mux.scala 19:72:@44117.4]
  wire [7:0] _T_97193; // @[Mux.scala 19:72:@44124.4]
  wire [15:0] _T_97201; // @[Mux.scala 19:72:@44132.4]
  wire [15:0] _T_97203; // @[Mux.scala 19:72:@44133.4]
  wire [7:0] _T_97210; // @[Mux.scala 19:72:@44140.4]
  wire [15:0] _T_97218; // @[Mux.scala 19:72:@44148.4]
  wire [15:0] _T_97220; // @[Mux.scala 19:72:@44149.4]
  wire [7:0] _T_97227; // @[Mux.scala 19:72:@44156.4]
  wire [15:0] _T_97235; // @[Mux.scala 19:72:@44164.4]
  wire [15:0] _T_97237; // @[Mux.scala 19:72:@44165.4]
  wire [7:0] _T_97244; // @[Mux.scala 19:72:@44172.4]
  wire [15:0] _T_97252; // @[Mux.scala 19:72:@44180.4]
  wire [15:0] _T_97254; // @[Mux.scala 19:72:@44181.4]
  wire [7:0] _T_97261; // @[Mux.scala 19:72:@44188.4]
  wire [15:0] _T_97269; // @[Mux.scala 19:72:@44196.4]
  wire [15:0] _T_97271; // @[Mux.scala 19:72:@44197.4]
  wire [7:0] _T_97278; // @[Mux.scala 19:72:@44204.4]
  wire [15:0] _T_97286; // @[Mux.scala 19:72:@44212.4]
  wire [15:0] _T_97288; // @[Mux.scala 19:72:@44213.4]
  wire [7:0] _T_97295; // @[Mux.scala 19:72:@44220.4]
  wire [15:0] _T_97303; // @[Mux.scala 19:72:@44228.4]
  wire [15:0] _T_97305; // @[Mux.scala 19:72:@44229.4]
  wire [7:0] _T_97312; // @[Mux.scala 19:72:@44236.4]
  wire [15:0] _T_97320; // @[Mux.scala 19:72:@44244.4]
  wire [15:0] _T_97322; // @[Mux.scala 19:72:@44245.4]
  wire [7:0] _T_97329; // @[Mux.scala 19:72:@44252.4]
  wire [15:0] _T_97337; // @[Mux.scala 19:72:@44260.4]
  wire [15:0] _T_97339; // @[Mux.scala 19:72:@44261.4]
  wire [7:0] _T_97346; // @[Mux.scala 19:72:@44268.4]
  wire [15:0] _T_97354; // @[Mux.scala 19:72:@44276.4]
  wire [15:0] _T_97356; // @[Mux.scala 19:72:@44277.4]
  wire [7:0] _T_97363; // @[Mux.scala 19:72:@44284.4]
  wire [15:0] _T_97371; // @[Mux.scala 19:72:@44292.4]
  wire [15:0] _T_97373; // @[Mux.scala 19:72:@44293.4]
  wire [7:0] _T_97380; // @[Mux.scala 19:72:@44300.4]
  wire [15:0] _T_97388; // @[Mux.scala 19:72:@44308.4]
  wire [15:0] _T_97390; // @[Mux.scala 19:72:@44309.4]
  wire [7:0] _T_97397; // @[Mux.scala 19:72:@44316.4]
  wire [15:0] _T_97405; // @[Mux.scala 19:72:@44324.4]
  wire [15:0] _T_97407; // @[Mux.scala 19:72:@44325.4]
  wire [15:0] _T_97408; // @[Mux.scala 19:72:@44326.4]
  wire [15:0] _T_97409; // @[Mux.scala 19:72:@44327.4]
  wire [15:0] _T_97410; // @[Mux.scala 19:72:@44328.4]
  wire [15:0] _T_97411; // @[Mux.scala 19:72:@44329.4]
  wire [15:0] _T_97412; // @[Mux.scala 19:72:@44330.4]
  wire [15:0] _T_97413; // @[Mux.scala 19:72:@44331.4]
  wire [15:0] _T_97414; // @[Mux.scala 19:72:@44332.4]
  wire [15:0] _T_97415; // @[Mux.scala 19:72:@44333.4]
  wire [15:0] _T_97416; // @[Mux.scala 19:72:@44334.4]
  wire [15:0] _T_97417; // @[Mux.scala 19:72:@44335.4]
  wire [15:0] _T_97418; // @[Mux.scala 19:72:@44336.4]
  wire [15:0] _T_97419; // @[Mux.scala 19:72:@44337.4]
  wire [15:0] _T_97420; // @[Mux.scala 19:72:@44338.4]
  wire [15:0] _T_97421; // @[Mux.scala 19:72:@44339.4]
  wire [15:0] _T_97422; // @[Mux.scala 19:72:@44340.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@44344.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@44346.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@44348.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@44350.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@44352.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@44354.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@44356.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@44358.4]
  wire  outputPriorityPorts_0_8; // @[Mux.scala 19:72:@44360.4]
  wire  outputPriorityPorts_0_9; // @[Mux.scala 19:72:@44362.4]
  wire  outputPriorityPorts_0_10; // @[Mux.scala 19:72:@44364.4]
  wire  outputPriorityPorts_0_11; // @[Mux.scala 19:72:@44366.4]
  wire  outputPriorityPorts_0_12; // @[Mux.scala 19:72:@44368.4]
  wire  outputPriorityPorts_0_13; // @[Mux.scala 19:72:@44370.4]
  wire  outputPriorityPorts_0_14; // @[Mux.scala 19:72:@44372.4]
  wire  outputPriorityPorts_0_15; // @[Mux.scala 19:72:@44374.4]
  wire  _T_97565; // @[LoadQueue.scala 313:47:@44396.6]
  wire [31:0] _GEN_2114; // @[LoadQueue.scala 314:36:@44400.6]
  wire  _GEN_2115; // @[LoadQueue.scala 314:36:@44400.6]
  wire  _GEN_2116; // @[LoadQueue.scala 308:34:@44392.4]
  wire [31:0] _GEN_2117; // @[LoadQueue.scala 308:34:@44392.4]
  wire  _T_97580; // @[LoadQueue.scala 313:47:@44409.6]
  wire [31:0] _GEN_2118; // @[LoadQueue.scala 314:36:@44413.6]
  wire  _GEN_2119; // @[LoadQueue.scala 314:36:@44413.6]
  wire  _GEN_2120; // @[LoadQueue.scala 308:34:@44405.4]
  wire [31:0] _GEN_2121; // @[LoadQueue.scala 308:34:@44405.4]
  wire  _T_97595; // @[LoadQueue.scala 313:47:@44422.6]
  wire [31:0] _GEN_2122; // @[LoadQueue.scala 314:36:@44426.6]
  wire  _GEN_2123; // @[LoadQueue.scala 314:36:@44426.6]
  wire  _GEN_2124; // @[LoadQueue.scala 308:34:@44418.4]
  wire [31:0] _GEN_2125; // @[LoadQueue.scala 308:34:@44418.4]
  wire  _T_97610; // @[LoadQueue.scala 313:47:@44435.6]
  wire [31:0] _GEN_2126; // @[LoadQueue.scala 314:36:@44439.6]
  wire  _GEN_2127; // @[LoadQueue.scala 314:36:@44439.6]
  wire  _GEN_2128; // @[LoadQueue.scala 308:34:@44431.4]
  wire [31:0] _GEN_2129; // @[LoadQueue.scala 308:34:@44431.4]
  wire  _T_97625; // @[LoadQueue.scala 313:47:@44448.6]
  wire [31:0] _GEN_2130; // @[LoadQueue.scala 314:36:@44452.6]
  wire  _GEN_2131; // @[LoadQueue.scala 314:36:@44452.6]
  wire  _GEN_2132; // @[LoadQueue.scala 308:34:@44444.4]
  wire [31:0] _GEN_2133; // @[LoadQueue.scala 308:34:@44444.4]
  wire  _T_97640; // @[LoadQueue.scala 313:47:@44461.6]
  wire [31:0] _GEN_2134; // @[LoadQueue.scala 314:36:@44465.6]
  wire  _GEN_2135; // @[LoadQueue.scala 314:36:@44465.6]
  wire  _GEN_2136; // @[LoadQueue.scala 308:34:@44457.4]
  wire [31:0] _GEN_2137; // @[LoadQueue.scala 308:34:@44457.4]
  wire  _T_97655; // @[LoadQueue.scala 313:47:@44474.6]
  wire [31:0] _GEN_2138; // @[LoadQueue.scala 314:36:@44478.6]
  wire  _GEN_2139; // @[LoadQueue.scala 314:36:@44478.6]
  wire  _GEN_2140; // @[LoadQueue.scala 308:34:@44470.4]
  wire [31:0] _GEN_2141; // @[LoadQueue.scala 308:34:@44470.4]
  wire  _T_97670; // @[LoadQueue.scala 313:47:@44487.6]
  wire [31:0] _GEN_2142; // @[LoadQueue.scala 314:36:@44491.6]
  wire  _GEN_2143; // @[LoadQueue.scala 314:36:@44491.6]
  wire  _GEN_2144; // @[LoadQueue.scala 308:34:@44483.4]
  wire [31:0] _GEN_2145; // @[LoadQueue.scala 308:34:@44483.4]
  wire  _T_97685; // @[LoadQueue.scala 313:47:@44500.6]
  wire [31:0] _GEN_2146; // @[LoadQueue.scala 314:36:@44504.6]
  wire  _GEN_2147; // @[LoadQueue.scala 314:36:@44504.6]
  wire  _GEN_2148; // @[LoadQueue.scala 308:34:@44496.4]
  wire [31:0] _GEN_2149; // @[LoadQueue.scala 308:34:@44496.4]
  wire  _T_97700; // @[LoadQueue.scala 313:47:@44513.6]
  wire [31:0] _GEN_2150; // @[LoadQueue.scala 314:36:@44517.6]
  wire  _GEN_2151; // @[LoadQueue.scala 314:36:@44517.6]
  wire  _GEN_2152; // @[LoadQueue.scala 308:34:@44509.4]
  wire [31:0] _GEN_2153; // @[LoadQueue.scala 308:34:@44509.4]
  wire  _T_97715; // @[LoadQueue.scala 313:47:@44526.6]
  wire [31:0] _GEN_2154; // @[LoadQueue.scala 314:36:@44530.6]
  wire  _GEN_2155; // @[LoadQueue.scala 314:36:@44530.6]
  wire  _GEN_2156; // @[LoadQueue.scala 308:34:@44522.4]
  wire [31:0] _GEN_2157; // @[LoadQueue.scala 308:34:@44522.4]
  wire  _T_97730; // @[LoadQueue.scala 313:47:@44539.6]
  wire [31:0] _GEN_2158; // @[LoadQueue.scala 314:36:@44543.6]
  wire  _GEN_2159; // @[LoadQueue.scala 314:36:@44543.6]
  wire  _GEN_2160; // @[LoadQueue.scala 308:34:@44535.4]
  wire [31:0] _GEN_2161; // @[LoadQueue.scala 308:34:@44535.4]
  wire  _T_97745; // @[LoadQueue.scala 313:47:@44552.6]
  wire [31:0] _GEN_2162; // @[LoadQueue.scala 314:36:@44556.6]
  wire  _GEN_2163; // @[LoadQueue.scala 314:36:@44556.6]
  wire  _GEN_2164; // @[LoadQueue.scala 308:34:@44548.4]
  wire [31:0] _GEN_2165; // @[LoadQueue.scala 308:34:@44548.4]
  wire  _T_97760; // @[LoadQueue.scala 313:47:@44565.6]
  wire [31:0] _GEN_2166; // @[LoadQueue.scala 314:36:@44569.6]
  wire  _GEN_2167; // @[LoadQueue.scala 314:36:@44569.6]
  wire  _GEN_2168; // @[LoadQueue.scala 308:34:@44561.4]
  wire [31:0] _GEN_2169; // @[LoadQueue.scala 308:34:@44561.4]
  wire  _T_97775; // @[LoadQueue.scala 313:47:@44578.6]
  wire [31:0] _GEN_2170; // @[LoadQueue.scala 314:36:@44582.6]
  wire  _GEN_2171; // @[LoadQueue.scala 314:36:@44582.6]
  wire  _GEN_2172; // @[LoadQueue.scala 308:34:@44574.4]
  wire [31:0] _GEN_2173; // @[LoadQueue.scala 308:34:@44574.4]
  wire  _T_97790; // @[LoadQueue.scala 313:47:@44591.6]
  wire [31:0] _GEN_2174; // @[LoadQueue.scala 314:36:@44595.6]
  wire  _GEN_2175; // @[LoadQueue.scala 314:36:@44595.6]
  wire  _GEN_2176; // @[LoadQueue.scala 308:34:@44587.4]
  wire [31:0] _GEN_2177; // @[LoadQueue.scala 308:34:@44587.4]
  wire  _T_97825; // @[LoadQueue.scala 326:108:@44601.4]
  wire  _T_97827; // @[LoadQueue.scala 327:34:@44602.4]
  wire  _T_97828; // @[LoadQueue.scala 327:31:@44603.4]
  wire  loadCompleting_0; // @[LoadQueue.scala 327:63:@44604.4]
  wire  _T_97839; // @[LoadQueue.scala 326:108:@44609.4]
  wire  _T_97841; // @[LoadQueue.scala 327:34:@44610.4]
  wire  _T_97842; // @[LoadQueue.scala 327:31:@44611.4]
  wire  loadCompleting_1; // @[LoadQueue.scala 327:63:@44612.4]
  wire  _T_97853; // @[LoadQueue.scala 326:108:@44617.4]
  wire  _T_97855; // @[LoadQueue.scala 327:34:@44618.4]
  wire  _T_97856; // @[LoadQueue.scala 327:31:@44619.4]
  wire  loadCompleting_2; // @[LoadQueue.scala 327:63:@44620.4]
  wire  _T_97867; // @[LoadQueue.scala 326:108:@44625.4]
  wire  _T_97869; // @[LoadQueue.scala 327:34:@44626.4]
  wire  _T_97870; // @[LoadQueue.scala 327:31:@44627.4]
  wire  loadCompleting_3; // @[LoadQueue.scala 327:63:@44628.4]
  wire  _T_97881; // @[LoadQueue.scala 326:108:@44633.4]
  wire  _T_97883; // @[LoadQueue.scala 327:34:@44634.4]
  wire  _T_97884; // @[LoadQueue.scala 327:31:@44635.4]
  wire  loadCompleting_4; // @[LoadQueue.scala 327:63:@44636.4]
  wire  _T_97895; // @[LoadQueue.scala 326:108:@44641.4]
  wire  _T_97897; // @[LoadQueue.scala 327:34:@44642.4]
  wire  _T_97898; // @[LoadQueue.scala 327:31:@44643.4]
  wire  loadCompleting_5; // @[LoadQueue.scala 327:63:@44644.4]
  wire  _T_97909; // @[LoadQueue.scala 326:108:@44649.4]
  wire  _T_97911; // @[LoadQueue.scala 327:34:@44650.4]
  wire  _T_97912; // @[LoadQueue.scala 327:31:@44651.4]
  wire  loadCompleting_6; // @[LoadQueue.scala 327:63:@44652.4]
  wire  _T_97923; // @[LoadQueue.scala 326:108:@44657.4]
  wire  _T_97925; // @[LoadQueue.scala 327:34:@44658.4]
  wire  _T_97926; // @[LoadQueue.scala 327:31:@44659.4]
  wire  loadCompleting_7; // @[LoadQueue.scala 327:63:@44660.4]
  wire  _T_97937; // @[LoadQueue.scala 326:108:@44665.4]
  wire  _T_97939; // @[LoadQueue.scala 327:34:@44666.4]
  wire  _T_97940; // @[LoadQueue.scala 327:31:@44667.4]
  wire  loadCompleting_8; // @[LoadQueue.scala 327:63:@44668.4]
  wire  _T_97951; // @[LoadQueue.scala 326:108:@44673.4]
  wire  _T_97953; // @[LoadQueue.scala 327:34:@44674.4]
  wire  _T_97954; // @[LoadQueue.scala 327:31:@44675.4]
  wire  loadCompleting_9; // @[LoadQueue.scala 327:63:@44676.4]
  wire  _T_97965; // @[LoadQueue.scala 326:108:@44681.4]
  wire  _T_97967; // @[LoadQueue.scala 327:34:@44682.4]
  wire  _T_97968; // @[LoadQueue.scala 327:31:@44683.4]
  wire  loadCompleting_10; // @[LoadQueue.scala 327:63:@44684.4]
  wire  _T_97979; // @[LoadQueue.scala 326:108:@44689.4]
  wire  _T_97981; // @[LoadQueue.scala 327:34:@44690.4]
  wire  _T_97982; // @[LoadQueue.scala 327:31:@44691.4]
  wire  loadCompleting_11; // @[LoadQueue.scala 327:63:@44692.4]
  wire  _T_97993; // @[LoadQueue.scala 326:108:@44697.4]
  wire  _T_97995; // @[LoadQueue.scala 327:34:@44698.4]
  wire  _T_97996; // @[LoadQueue.scala 327:31:@44699.4]
  wire  loadCompleting_12; // @[LoadQueue.scala 327:63:@44700.4]
  wire  _T_98007; // @[LoadQueue.scala 326:108:@44705.4]
  wire  _T_98009; // @[LoadQueue.scala 327:34:@44706.4]
  wire  _T_98010; // @[LoadQueue.scala 327:31:@44707.4]
  wire  loadCompleting_13; // @[LoadQueue.scala 327:63:@44708.4]
  wire  _T_98021; // @[LoadQueue.scala 326:108:@44713.4]
  wire  _T_98023; // @[LoadQueue.scala 327:34:@44714.4]
  wire  _T_98024; // @[LoadQueue.scala 327:31:@44715.4]
  wire  loadCompleting_14; // @[LoadQueue.scala 327:63:@44716.4]
  wire  _T_98035; // @[LoadQueue.scala 326:108:@44721.4]
  wire  _T_98037; // @[LoadQueue.scala 327:34:@44722.4]
  wire  _T_98038; // @[LoadQueue.scala 327:31:@44723.4]
  wire  loadCompleting_15; // @[LoadQueue.scala 327:63:@44724.4]
  wire  _GEN_2178; // @[LoadQueue.scala 337:46:@44733.6]
  wire  _GEN_2179; // @[LoadQueue.scala 335:34:@44729.4]
  wire  _GEN_2180; // @[LoadQueue.scala 337:46:@44740.6]
  wire  _GEN_2181; // @[LoadQueue.scala 335:34:@44736.4]
  wire  _GEN_2182; // @[LoadQueue.scala 337:46:@44747.6]
  wire  _GEN_2183; // @[LoadQueue.scala 335:34:@44743.4]
  wire  _GEN_2184; // @[LoadQueue.scala 337:46:@44754.6]
  wire  _GEN_2185; // @[LoadQueue.scala 335:34:@44750.4]
  wire  _GEN_2186; // @[LoadQueue.scala 337:46:@44761.6]
  wire  _GEN_2187; // @[LoadQueue.scala 335:34:@44757.4]
  wire  _GEN_2188; // @[LoadQueue.scala 337:46:@44768.6]
  wire  _GEN_2189; // @[LoadQueue.scala 335:34:@44764.4]
  wire  _GEN_2190; // @[LoadQueue.scala 337:46:@44775.6]
  wire  _GEN_2191; // @[LoadQueue.scala 335:34:@44771.4]
  wire  _GEN_2192; // @[LoadQueue.scala 337:46:@44782.6]
  wire  _GEN_2193; // @[LoadQueue.scala 335:34:@44778.4]
  wire  _GEN_2194; // @[LoadQueue.scala 337:46:@44789.6]
  wire  _GEN_2195; // @[LoadQueue.scala 335:34:@44785.4]
  wire  _GEN_2196; // @[LoadQueue.scala 337:46:@44796.6]
  wire  _GEN_2197; // @[LoadQueue.scala 335:34:@44792.4]
  wire  _GEN_2198; // @[LoadQueue.scala 337:46:@44803.6]
  wire  _GEN_2199; // @[LoadQueue.scala 335:34:@44799.4]
  wire  _GEN_2200; // @[LoadQueue.scala 337:46:@44810.6]
  wire  _GEN_2201; // @[LoadQueue.scala 335:34:@44806.4]
  wire  _GEN_2202; // @[LoadQueue.scala 337:46:@44817.6]
  wire  _GEN_2203; // @[LoadQueue.scala 335:34:@44813.4]
  wire  _GEN_2204; // @[LoadQueue.scala 337:46:@44824.6]
  wire  _GEN_2205; // @[LoadQueue.scala 335:34:@44820.4]
  wire  _GEN_2206; // @[LoadQueue.scala 337:46:@44831.6]
  wire  _GEN_2207; // @[LoadQueue.scala 335:34:@44827.4]
  wire  _GEN_2208; // @[LoadQueue.scala 337:46:@44838.6]
  wire  _GEN_2209; // @[LoadQueue.scala 335:34:@44834.4]
  wire  _T_98169; // @[LoadQueue.scala 348:24:@44907.4]
  wire  _T_98170; // @[LoadQueue.scala 348:24:@44908.4]
  wire  _T_98171; // @[LoadQueue.scala 348:24:@44909.4]
  wire  _T_98172; // @[LoadQueue.scala 348:24:@44910.4]
  wire  _T_98173; // @[LoadQueue.scala 348:24:@44911.4]
  wire  _T_98174; // @[LoadQueue.scala 348:24:@44912.4]
  wire  _T_98175; // @[LoadQueue.scala 348:24:@44913.4]
  wire  _T_98176; // @[LoadQueue.scala 348:24:@44914.4]
  wire  _T_98177; // @[LoadQueue.scala 348:24:@44915.4]
  wire  _T_98178; // @[LoadQueue.scala 348:24:@44916.4]
  wire  _T_98179; // @[LoadQueue.scala 348:24:@44917.4]
  wire  _T_98180; // @[LoadQueue.scala 348:24:@44918.4]
  wire  _T_98181; // @[LoadQueue.scala 348:24:@44919.4]
  wire  _T_98182; // @[LoadQueue.scala 348:24:@44920.4]
  wire  _T_98183; // @[LoadQueue.scala 348:24:@44921.4]
  wire [3:0] _T_98200; // @[Mux.scala 31:69:@44923.6]
  wire [3:0] _T_98201; // @[Mux.scala 31:69:@44924.6]
  wire [3:0] _T_98202; // @[Mux.scala 31:69:@44925.6]
  wire [3:0] _T_98203; // @[Mux.scala 31:69:@44926.6]
  wire [3:0] _T_98204; // @[Mux.scala 31:69:@44927.6]
  wire [3:0] _T_98205; // @[Mux.scala 31:69:@44928.6]
  wire [3:0] _T_98206; // @[Mux.scala 31:69:@44929.6]
  wire [3:0] _T_98207; // @[Mux.scala 31:69:@44930.6]
  wire [3:0] _T_98208; // @[Mux.scala 31:69:@44931.6]
  wire [3:0] _T_98209; // @[Mux.scala 31:69:@44932.6]
  wire [3:0] _T_98210; // @[Mux.scala 31:69:@44933.6]
  wire [3:0] _T_98211; // @[Mux.scala 31:69:@44934.6]
  wire [3:0] _T_98212; // @[Mux.scala 31:69:@44935.6]
  wire [3:0] _T_98213; // @[Mux.scala 31:69:@44936.6]
  wire [3:0] _T_98214; // @[Mux.scala 31:69:@44937.6]
  wire [31:0] _GEN_2211; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2212; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2213; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2214; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2215; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2216; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2217; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2218; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2219; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2220; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2221; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2222; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2223; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2224; // @[LoadQueue.scala 349:37:@44938.6]
  wire [31:0] _GEN_2225; // @[LoadQueue.scala 349:37:@44938.6]
  wire  _GEN_2229; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2230; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2231; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2232; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2233; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2234; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2235; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2236; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2237; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2238; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2239; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2240; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2241; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2242; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2243; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2245; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2246; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2247; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2248; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2249; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2250; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2251; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2252; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2253; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2254; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2255; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2256; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2257; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2258; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _GEN_2259; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _T_98225; // @[LoadQueue.scala 363:29:@44945.4]
  wire  _T_98226; // @[LoadQueue.scala 363:63:@44946.4]
  wire  _T_98228; // @[LoadQueue.scala 363:75:@44947.4]
  wire  _T_98229; // @[LoadQueue.scala 363:72:@44948.4]
  wire  _T_98230; // @[LoadQueue.scala 363:54:@44949.4]
  wire [4:0] _T_98233; // @[util.scala 10:8:@44951.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@44952.6]
  wire [4:0] _T_98234; // @[util.scala 10:14:@44952.6]
  wire [4:0] _GEN_2260; // @[LoadQueue.scala 363:91:@44950.4]
  wire [3:0] _GEN_2358; // @[util.scala 10:8:@44956.6]
  wire [4:0] _T_98236; // @[util.scala 10:8:@44956.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@44957.6]
  wire [4:0] _T_98237; // @[util.scala 10:14:@44957.6]
  wire [4:0] _GEN_2261; // @[LoadQueue.scala 367:20:@44955.4]
  wire  _T_98239; // @[LoadQueue.scala 371:82:@44960.4]
  wire  _T_98240; // @[LoadQueue.scala 371:79:@44961.4]
  wire  _T_98242; // @[LoadQueue.scala 371:82:@44962.4]
  wire  _T_98243; // @[LoadQueue.scala 371:79:@44963.4]
  wire  _T_98245; // @[LoadQueue.scala 371:82:@44964.4]
  wire  _T_98246; // @[LoadQueue.scala 371:79:@44965.4]
  wire  _T_98248; // @[LoadQueue.scala 371:82:@44966.4]
  wire  _T_98249; // @[LoadQueue.scala 371:79:@44967.4]
  wire  _T_98251; // @[LoadQueue.scala 371:82:@44968.4]
  wire  _T_98252; // @[LoadQueue.scala 371:79:@44969.4]
  wire  _T_98254; // @[LoadQueue.scala 371:82:@44970.4]
  wire  _T_98255; // @[LoadQueue.scala 371:79:@44971.4]
  wire  _T_98257; // @[LoadQueue.scala 371:82:@44972.4]
  wire  _T_98258; // @[LoadQueue.scala 371:79:@44973.4]
  wire  _T_98260; // @[LoadQueue.scala 371:82:@44974.4]
  wire  _T_98261; // @[LoadQueue.scala 371:79:@44975.4]
  wire  _T_98263; // @[LoadQueue.scala 371:82:@44976.4]
  wire  _T_98264; // @[LoadQueue.scala 371:79:@44977.4]
  wire  _T_98266; // @[LoadQueue.scala 371:82:@44978.4]
  wire  _T_98267; // @[LoadQueue.scala 371:79:@44979.4]
  wire  _T_98269; // @[LoadQueue.scala 371:82:@44980.4]
  wire  _T_98270; // @[LoadQueue.scala 371:79:@44981.4]
  wire  _T_98272; // @[LoadQueue.scala 371:82:@44982.4]
  wire  _T_98273; // @[LoadQueue.scala 371:79:@44983.4]
  wire  _T_98275; // @[LoadQueue.scala 371:82:@44984.4]
  wire  _T_98276; // @[LoadQueue.scala 371:79:@44985.4]
  wire  _T_98278; // @[LoadQueue.scala 371:82:@44986.4]
  wire  _T_98279; // @[LoadQueue.scala 371:79:@44987.4]
  wire  _T_98281; // @[LoadQueue.scala 371:82:@44988.4]
  wire  _T_98282; // @[LoadQueue.scala 371:79:@44989.4]
  wire  _T_98284; // @[LoadQueue.scala 371:82:@44990.4]
  wire  _T_98285; // @[LoadQueue.scala 371:79:@44991.4]
  wire  _T_98310; // @[LoadQueue.scala 371:96:@45010.4]
  wire  _T_98311; // @[LoadQueue.scala 371:96:@45011.4]
  wire  _T_98312; // @[LoadQueue.scala 371:96:@45012.4]
  wire  _T_98313; // @[LoadQueue.scala 371:96:@45013.4]
  wire  _T_98314; // @[LoadQueue.scala 371:96:@45014.4]
  wire  _T_98315; // @[LoadQueue.scala 371:96:@45015.4]
  wire  _T_98316; // @[LoadQueue.scala 371:96:@45016.4]
  wire  _T_98317; // @[LoadQueue.scala 371:96:@45017.4]
  wire  _T_98318; // @[LoadQueue.scala 371:96:@45018.4]
  wire  _T_98319; // @[LoadQueue.scala 371:96:@45019.4]
  wire  _T_98320; // @[LoadQueue.scala 371:96:@45020.4]
  wire  _T_98321; // @[LoadQueue.scala 371:96:@45021.4]
  wire  _T_98322; // @[LoadQueue.scala 371:96:@45022.4]
  wire  _T_98323; // @[LoadQueue.scala 371:96:@45023.4]
  assign _GEN_2262 = {{2'd0}, tail}; // @[util.scala 14:20:@7670.4]
  assign _T_1716 = 6'h10 - _GEN_2262; // @[util.scala 14:20:@7670.4]
  assign _T_1717 = $unsigned(_T_1716); // @[util.scala 14:20:@7671.4]
  assign _T_1718 = _T_1717[5:0]; // @[util.scala 14:20:@7672.4]
  assign _GEN_0 = _T_1718 % 6'h10; // @[util.scala 14:25:@7673.4]
  assign _T_1719 = _GEN_0[4:0]; // @[util.scala 14:25:@7673.4]
  assign _GEN_2263 = {{4'd0}, io_bbNumLoads}; // @[LoadQueue.scala 71:46:@7674.4]
  assign _T_1720 = _T_1719 < _GEN_2263; // @[LoadQueue.scala 71:46:@7674.4]
  assign initBits_0 = _T_1720 & io_bbStart; // @[LoadQueue.scala 71:63:@7675.4]
  assign _T_1725 = 6'h11 - _GEN_2262; // @[util.scala 14:20:@7677.4]
  assign _T_1726 = $unsigned(_T_1725); // @[util.scala 14:20:@7678.4]
  assign _T_1727 = _T_1726[5:0]; // @[util.scala 14:20:@7679.4]
  assign _GEN_16 = _T_1727 % 6'h10; // @[util.scala 14:25:@7680.4]
  assign _T_1728 = _GEN_16[4:0]; // @[util.scala 14:25:@7680.4]
  assign _T_1729 = _T_1728 < _GEN_2263; // @[LoadQueue.scala 71:46:@7681.4]
  assign initBits_1 = _T_1729 & io_bbStart; // @[LoadQueue.scala 71:63:@7682.4]
  assign _T_1734 = 6'h12 - _GEN_2262; // @[util.scala 14:20:@7684.4]
  assign _T_1735 = $unsigned(_T_1734); // @[util.scala 14:20:@7685.4]
  assign _T_1736 = _T_1735[5:0]; // @[util.scala 14:20:@7686.4]
  assign _GEN_17 = _T_1736 % 6'h10; // @[util.scala 14:25:@7687.4]
  assign _T_1737 = _GEN_17[4:0]; // @[util.scala 14:25:@7687.4]
  assign _T_1738 = _T_1737 < _GEN_2263; // @[LoadQueue.scala 71:46:@7688.4]
  assign initBits_2 = _T_1738 & io_bbStart; // @[LoadQueue.scala 71:63:@7689.4]
  assign _T_1743 = 6'h13 - _GEN_2262; // @[util.scala 14:20:@7691.4]
  assign _T_1744 = $unsigned(_T_1743); // @[util.scala 14:20:@7692.4]
  assign _T_1745 = _T_1744[5:0]; // @[util.scala 14:20:@7693.4]
  assign _GEN_18 = _T_1745 % 6'h10; // @[util.scala 14:25:@7694.4]
  assign _T_1746 = _GEN_18[4:0]; // @[util.scala 14:25:@7694.4]
  assign _T_1747 = _T_1746 < _GEN_2263; // @[LoadQueue.scala 71:46:@7695.4]
  assign initBits_3 = _T_1747 & io_bbStart; // @[LoadQueue.scala 71:63:@7696.4]
  assign _T_1752 = 6'h14 - _GEN_2262; // @[util.scala 14:20:@7698.4]
  assign _T_1753 = $unsigned(_T_1752); // @[util.scala 14:20:@7699.4]
  assign _T_1754 = _T_1753[5:0]; // @[util.scala 14:20:@7700.4]
  assign _GEN_19 = _T_1754 % 6'h10; // @[util.scala 14:25:@7701.4]
  assign _T_1755 = _GEN_19[4:0]; // @[util.scala 14:25:@7701.4]
  assign _T_1756 = _T_1755 < _GEN_2263; // @[LoadQueue.scala 71:46:@7702.4]
  assign initBits_4 = _T_1756 & io_bbStart; // @[LoadQueue.scala 71:63:@7703.4]
  assign _T_1761 = 6'h15 - _GEN_2262; // @[util.scala 14:20:@7705.4]
  assign _T_1762 = $unsigned(_T_1761); // @[util.scala 14:20:@7706.4]
  assign _T_1763 = _T_1762[5:0]; // @[util.scala 14:20:@7707.4]
  assign _GEN_20 = _T_1763 % 6'h10; // @[util.scala 14:25:@7708.4]
  assign _T_1764 = _GEN_20[4:0]; // @[util.scala 14:25:@7708.4]
  assign _T_1765 = _T_1764 < _GEN_2263; // @[LoadQueue.scala 71:46:@7709.4]
  assign initBits_5 = _T_1765 & io_bbStart; // @[LoadQueue.scala 71:63:@7710.4]
  assign _T_1770 = 6'h16 - _GEN_2262; // @[util.scala 14:20:@7712.4]
  assign _T_1771 = $unsigned(_T_1770); // @[util.scala 14:20:@7713.4]
  assign _T_1772 = _T_1771[5:0]; // @[util.scala 14:20:@7714.4]
  assign _GEN_21 = _T_1772 % 6'h10; // @[util.scala 14:25:@7715.4]
  assign _T_1773 = _GEN_21[4:0]; // @[util.scala 14:25:@7715.4]
  assign _T_1774 = _T_1773 < _GEN_2263; // @[LoadQueue.scala 71:46:@7716.4]
  assign initBits_6 = _T_1774 & io_bbStart; // @[LoadQueue.scala 71:63:@7717.4]
  assign _T_1779 = 6'h17 - _GEN_2262; // @[util.scala 14:20:@7719.4]
  assign _T_1780 = $unsigned(_T_1779); // @[util.scala 14:20:@7720.4]
  assign _T_1781 = _T_1780[5:0]; // @[util.scala 14:20:@7721.4]
  assign _GEN_22 = _T_1781 % 6'h10; // @[util.scala 14:25:@7722.4]
  assign _T_1782 = _GEN_22[4:0]; // @[util.scala 14:25:@7722.4]
  assign _T_1783 = _T_1782 < _GEN_2263; // @[LoadQueue.scala 71:46:@7723.4]
  assign initBits_7 = _T_1783 & io_bbStart; // @[LoadQueue.scala 71:63:@7724.4]
  assign _T_1788 = 6'h18 - _GEN_2262; // @[util.scala 14:20:@7726.4]
  assign _T_1789 = $unsigned(_T_1788); // @[util.scala 14:20:@7727.4]
  assign _T_1790 = _T_1789[5:0]; // @[util.scala 14:20:@7728.4]
  assign _GEN_23 = _T_1790 % 6'h10; // @[util.scala 14:25:@7729.4]
  assign _T_1791 = _GEN_23[4:0]; // @[util.scala 14:25:@7729.4]
  assign _T_1792 = _T_1791 < _GEN_2263; // @[LoadQueue.scala 71:46:@7730.4]
  assign initBits_8 = _T_1792 & io_bbStart; // @[LoadQueue.scala 71:63:@7731.4]
  assign _T_1797 = 6'h19 - _GEN_2262; // @[util.scala 14:20:@7733.4]
  assign _T_1798 = $unsigned(_T_1797); // @[util.scala 14:20:@7734.4]
  assign _T_1799 = _T_1798[5:0]; // @[util.scala 14:20:@7735.4]
  assign _GEN_24 = _T_1799 % 6'h10; // @[util.scala 14:25:@7736.4]
  assign _T_1800 = _GEN_24[4:0]; // @[util.scala 14:25:@7736.4]
  assign _T_1801 = _T_1800 < _GEN_2263; // @[LoadQueue.scala 71:46:@7737.4]
  assign initBits_9 = _T_1801 & io_bbStart; // @[LoadQueue.scala 71:63:@7738.4]
  assign _T_1806 = 6'h1a - _GEN_2262; // @[util.scala 14:20:@7740.4]
  assign _T_1807 = $unsigned(_T_1806); // @[util.scala 14:20:@7741.4]
  assign _T_1808 = _T_1807[5:0]; // @[util.scala 14:20:@7742.4]
  assign _GEN_25 = _T_1808 % 6'h10; // @[util.scala 14:25:@7743.4]
  assign _T_1809 = _GEN_25[4:0]; // @[util.scala 14:25:@7743.4]
  assign _T_1810 = _T_1809 < _GEN_2263; // @[LoadQueue.scala 71:46:@7744.4]
  assign initBits_10 = _T_1810 & io_bbStart; // @[LoadQueue.scala 71:63:@7745.4]
  assign _T_1815 = 6'h1b - _GEN_2262; // @[util.scala 14:20:@7747.4]
  assign _T_1816 = $unsigned(_T_1815); // @[util.scala 14:20:@7748.4]
  assign _T_1817 = _T_1816[5:0]; // @[util.scala 14:20:@7749.4]
  assign _GEN_26 = _T_1817 % 6'h10; // @[util.scala 14:25:@7750.4]
  assign _T_1818 = _GEN_26[4:0]; // @[util.scala 14:25:@7750.4]
  assign _T_1819 = _T_1818 < _GEN_2263; // @[LoadQueue.scala 71:46:@7751.4]
  assign initBits_11 = _T_1819 & io_bbStart; // @[LoadQueue.scala 71:63:@7752.4]
  assign _T_1824 = 6'h1c - _GEN_2262; // @[util.scala 14:20:@7754.4]
  assign _T_1825 = $unsigned(_T_1824); // @[util.scala 14:20:@7755.4]
  assign _T_1826 = _T_1825[5:0]; // @[util.scala 14:20:@7756.4]
  assign _GEN_27 = _T_1826 % 6'h10; // @[util.scala 14:25:@7757.4]
  assign _T_1827 = _GEN_27[4:0]; // @[util.scala 14:25:@7757.4]
  assign _T_1828 = _T_1827 < _GEN_2263; // @[LoadQueue.scala 71:46:@7758.4]
  assign initBits_12 = _T_1828 & io_bbStart; // @[LoadQueue.scala 71:63:@7759.4]
  assign _T_1833 = 6'h1d - _GEN_2262; // @[util.scala 14:20:@7761.4]
  assign _T_1834 = $unsigned(_T_1833); // @[util.scala 14:20:@7762.4]
  assign _T_1835 = _T_1834[5:0]; // @[util.scala 14:20:@7763.4]
  assign _GEN_28 = _T_1835 % 6'h10; // @[util.scala 14:25:@7764.4]
  assign _T_1836 = _GEN_28[4:0]; // @[util.scala 14:25:@7764.4]
  assign _T_1837 = _T_1836 < _GEN_2263; // @[LoadQueue.scala 71:46:@7765.4]
  assign initBits_13 = _T_1837 & io_bbStart; // @[LoadQueue.scala 71:63:@7766.4]
  assign _T_1842 = 6'h1e - _GEN_2262; // @[util.scala 14:20:@7768.4]
  assign _T_1843 = $unsigned(_T_1842); // @[util.scala 14:20:@7769.4]
  assign _T_1844 = _T_1843[5:0]; // @[util.scala 14:20:@7770.4]
  assign _GEN_29 = _T_1844 % 6'h10; // @[util.scala 14:25:@7771.4]
  assign _T_1845 = _GEN_29[4:0]; // @[util.scala 14:25:@7771.4]
  assign _T_1846 = _T_1845 < _GEN_2263; // @[LoadQueue.scala 71:46:@7772.4]
  assign initBits_14 = _T_1846 & io_bbStart; // @[LoadQueue.scala 71:63:@7773.4]
  assign _T_1851 = 6'h1f - _GEN_2262; // @[util.scala 14:20:@7775.4]
  assign _T_1852 = $unsigned(_T_1851); // @[util.scala 14:20:@7776.4]
  assign _T_1853 = _T_1852[5:0]; // @[util.scala 14:20:@7777.4]
  assign _GEN_30 = _T_1853 % 6'h10; // @[util.scala 14:25:@7778.4]
  assign _T_1854 = _GEN_30[4:0]; // @[util.scala 14:25:@7778.4]
  assign _T_1855 = _T_1854 < _GEN_2263; // @[LoadQueue.scala 71:46:@7779.4]
  assign initBits_15 = _T_1855 & io_bbStart; // @[LoadQueue.scala 71:63:@7780.4]
  assign _T_1878 = allocatedEntries_0 | initBits_0; // @[LoadQueue.scala 73:78:@7798.4]
  assign _T_1879 = allocatedEntries_1 | initBits_1; // @[LoadQueue.scala 73:78:@7799.4]
  assign _T_1880 = allocatedEntries_2 | initBits_2; // @[LoadQueue.scala 73:78:@7800.4]
  assign _T_1881 = allocatedEntries_3 | initBits_3; // @[LoadQueue.scala 73:78:@7801.4]
  assign _T_1882 = allocatedEntries_4 | initBits_4; // @[LoadQueue.scala 73:78:@7802.4]
  assign _T_1883 = allocatedEntries_5 | initBits_5; // @[LoadQueue.scala 73:78:@7803.4]
  assign _T_1884 = allocatedEntries_6 | initBits_6; // @[LoadQueue.scala 73:78:@7804.4]
  assign _T_1885 = allocatedEntries_7 | initBits_7; // @[LoadQueue.scala 73:78:@7805.4]
  assign _T_1886 = allocatedEntries_8 | initBits_8; // @[LoadQueue.scala 73:78:@7806.4]
  assign _T_1887 = allocatedEntries_9 | initBits_9; // @[LoadQueue.scala 73:78:@7807.4]
  assign _T_1888 = allocatedEntries_10 | initBits_10; // @[LoadQueue.scala 73:78:@7808.4]
  assign _T_1889 = allocatedEntries_11 | initBits_11; // @[LoadQueue.scala 73:78:@7809.4]
  assign _T_1890 = allocatedEntries_12 | initBits_12; // @[LoadQueue.scala 73:78:@7810.4]
  assign _T_1891 = allocatedEntries_13 | initBits_13; // @[LoadQueue.scala 73:78:@7811.4]
  assign _T_1892 = allocatedEntries_14 | initBits_14; // @[LoadQueue.scala 73:78:@7812.4]
  assign _T_1893 = allocatedEntries_15 | initBits_15; // @[LoadQueue.scala 73:78:@7813.4]
  assign _T_1924 = _T_1719[3:0]; // @[:@7853.6]
  assign _GEN_1 = 4'h1 == _T_1924 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_2 = 4'h2 == _T_1924 ? io_bbLoadOffsets_2 : _GEN_1; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_3 = 4'h3 == _T_1924 ? io_bbLoadOffsets_3 : _GEN_2; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_4 = 4'h4 == _T_1924 ? io_bbLoadOffsets_4 : _GEN_3; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_5 = 4'h5 == _T_1924 ? io_bbLoadOffsets_5 : _GEN_4; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_6 = 4'h6 == _T_1924 ? io_bbLoadOffsets_6 : _GEN_5; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_7 = 4'h7 == _T_1924 ? io_bbLoadOffsets_7 : _GEN_6; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_8 = 4'h8 == _T_1924 ? io_bbLoadOffsets_8 : _GEN_7; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_9 = 4'h9 == _T_1924 ? io_bbLoadOffsets_9 : _GEN_8; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_10 = 4'ha == _T_1924 ? io_bbLoadOffsets_10 : _GEN_9; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_11 = 4'hb == _T_1924 ? io_bbLoadOffsets_11 : _GEN_10; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_12 = 4'hc == _T_1924 ? io_bbLoadOffsets_12 : _GEN_11; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_13 = 4'hd == _T_1924 ? io_bbLoadOffsets_13 : _GEN_12; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_14 = 4'he == _T_1924 ? io_bbLoadOffsets_14 : _GEN_13; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_15 = 4'hf == _T_1924 ? io_bbLoadOffsets_15 : _GEN_14; // @[LoadQueue.scala 77:20:@7854.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[LoadQueue.scala 76:25:@7847.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[LoadQueue.scala 76:25:@7847.4]
  assign _T_1942 = _T_1728[3:0]; // @[:@7869.6]
  assign _GEN_35 = 4'h1 == _T_1942 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_36 = 4'h2 == _T_1942 ? io_bbLoadOffsets_2 : _GEN_35; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_37 = 4'h3 == _T_1942 ? io_bbLoadOffsets_3 : _GEN_36; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_38 = 4'h4 == _T_1942 ? io_bbLoadOffsets_4 : _GEN_37; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_39 = 4'h5 == _T_1942 ? io_bbLoadOffsets_5 : _GEN_38; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_40 = 4'h6 == _T_1942 ? io_bbLoadOffsets_6 : _GEN_39; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_41 = 4'h7 == _T_1942 ? io_bbLoadOffsets_7 : _GEN_40; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_42 = 4'h8 == _T_1942 ? io_bbLoadOffsets_8 : _GEN_41; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_43 = 4'h9 == _T_1942 ? io_bbLoadOffsets_9 : _GEN_42; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_44 = 4'ha == _T_1942 ? io_bbLoadOffsets_10 : _GEN_43; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_45 = 4'hb == _T_1942 ? io_bbLoadOffsets_11 : _GEN_44; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_46 = 4'hc == _T_1942 ? io_bbLoadOffsets_12 : _GEN_45; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_47 = 4'hd == _T_1942 ? io_bbLoadOffsets_13 : _GEN_46; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_48 = 4'he == _T_1942 ? io_bbLoadOffsets_14 : _GEN_47; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_49 = 4'hf == _T_1942 ? io_bbLoadOffsets_15 : _GEN_48; // @[LoadQueue.scala 77:20:@7870.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[LoadQueue.scala 76:25:@7863.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[LoadQueue.scala 76:25:@7863.4]
  assign _T_1960 = _T_1737[3:0]; // @[:@7885.6]
  assign _GEN_69 = 4'h1 == _T_1960 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_70 = 4'h2 == _T_1960 ? io_bbLoadOffsets_2 : _GEN_69; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_71 = 4'h3 == _T_1960 ? io_bbLoadOffsets_3 : _GEN_70; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_72 = 4'h4 == _T_1960 ? io_bbLoadOffsets_4 : _GEN_71; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_73 = 4'h5 == _T_1960 ? io_bbLoadOffsets_5 : _GEN_72; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_74 = 4'h6 == _T_1960 ? io_bbLoadOffsets_6 : _GEN_73; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_75 = 4'h7 == _T_1960 ? io_bbLoadOffsets_7 : _GEN_74; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_76 = 4'h8 == _T_1960 ? io_bbLoadOffsets_8 : _GEN_75; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_77 = 4'h9 == _T_1960 ? io_bbLoadOffsets_9 : _GEN_76; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_78 = 4'ha == _T_1960 ? io_bbLoadOffsets_10 : _GEN_77; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_79 = 4'hb == _T_1960 ? io_bbLoadOffsets_11 : _GEN_78; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_80 = 4'hc == _T_1960 ? io_bbLoadOffsets_12 : _GEN_79; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_81 = 4'hd == _T_1960 ? io_bbLoadOffsets_13 : _GEN_80; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_82 = 4'he == _T_1960 ? io_bbLoadOffsets_14 : _GEN_81; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_83 = 4'hf == _T_1960 ? io_bbLoadOffsets_15 : _GEN_82; // @[LoadQueue.scala 77:20:@7886.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[LoadQueue.scala 76:25:@7879.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[LoadQueue.scala 76:25:@7879.4]
  assign _T_1978 = _T_1746[3:0]; // @[:@7901.6]
  assign _GEN_103 = 4'h1 == _T_1978 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_104 = 4'h2 == _T_1978 ? io_bbLoadOffsets_2 : _GEN_103; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_105 = 4'h3 == _T_1978 ? io_bbLoadOffsets_3 : _GEN_104; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_106 = 4'h4 == _T_1978 ? io_bbLoadOffsets_4 : _GEN_105; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_107 = 4'h5 == _T_1978 ? io_bbLoadOffsets_5 : _GEN_106; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_108 = 4'h6 == _T_1978 ? io_bbLoadOffsets_6 : _GEN_107; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_109 = 4'h7 == _T_1978 ? io_bbLoadOffsets_7 : _GEN_108; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_110 = 4'h8 == _T_1978 ? io_bbLoadOffsets_8 : _GEN_109; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_111 = 4'h9 == _T_1978 ? io_bbLoadOffsets_9 : _GEN_110; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_112 = 4'ha == _T_1978 ? io_bbLoadOffsets_10 : _GEN_111; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_113 = 4'hb == _T_1978 ? io_bbLoadOffsets_11 : _GEN_112; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_114 = 4'hc == _T_1978 ? io_bbLoadOffsets_12 : _GEN_113; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_115 = 4'hd == _T_1978 ? io_bbLoadOffsets_13 : _GEN_114; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_116 = 4'he == _T_1978 ? io_bbLoadOffsets_14 : _GEN_115; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_117 = 4'hf == _T_1978 ? io_bbLoadOffsets_15 : _GEN_116; // @[LoadQueue.scala 77:20:@7902.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[LoadQueue.scala 76:25:@7895.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[LoadQueue.scala 76:25:@7895.4]
  assign _T_1996 = _T_1755[3:0]; // @[:@7917.6]
  assign _GEN_137 = 4'h1 == _T_1996 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_138 = 4'h2 == _T_1996 ? io_bbLoadOffsets_2 : _GEN_137; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_139 = 4'h3 == _T_1996 ? io_bbLoadOffsets_3 : _GEN_138; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_140 = 4'h4 == _T_1996 ? io_bbLoadOffsets_4 : _GEN_139; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_141 = 4'h5 == _T_1996 ? io_bbLoadOffsets_5 : _GEN_140; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_142 = 4'h6 == _T_1996 ? io_bbLoadOffsets_6 : _GEN_141; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_143 = 4'h7 == _T_1996 ? io_bbLoadOffsets_7 : _GEN_142; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_144 = 4'h8 == _T_1996 ? io_bbLoadOffsets_8 : _GEN_143; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_145 = 4'h9 == _T_1996 ? io_bbLoadOffsets_9 : _GEN_144; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_146 = 4'ha == _T_1996 ? io_bbLoadOffsets_10 : _GEN_145; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_147 = 4'hb == _T_1996 ? io_bbLoadOffsets_11 : _GEN_146; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_148 = 4'hc == _T_1996 ? io_bbLoadOffsets_12 : _GEN_147; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_149 = 4'hd == _T_1996 ? io_bbLoadOffsets_13 : _GEN_148; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_150 = 4'he == _T_1996 ? io_bbLoadOffsets_14 : _GEN_149; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_151 = 4'hf == _T_1996 ? io_bbLoadOffsets_15 : _GEN_150; // @[LoadQueue.scala 77:20:@7918.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[LoadQueue.scala 76:25:@7911.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[LoadQueue.scala 76:25:@7911.4]
  assign _T_2014 = _T_1764[3:0]; // @[:@7933.6]
  assign _GEN_171 = 4'h1 == _T_2014 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_172 = 4'h2 == _T_2014 ? io_bbLoadOffsets_2 : _GEN_171; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_173 = 4'h3 == _T_2014 ? io_bbLoadOffsets_3 : _GEN_172; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_174 = 4'h4 == _T_2014 ? io_bbLoadOffsets_4 : _GEN_173; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_175 = 4'h5 == _T_2014 ? io_bbLoadOffsets_5 : _GEN_174; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_176 = 4'h6 == _T_2014 ? io_bbLoadOffsets_6 : _GEN_175; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_177 = 4'h7 == _T_2014 ? io_bbLoadOffsets_7 : _GEN_176; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_178 = 4'h8 == _T_2014 ? io_bbLoadOffsets_8 : _GEN_177; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_179 = 4'h9 == _T_2014 ? io_bbLoadOffsets_9 : _GEN_178; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_180 = 4'ha == _T_2014 ? io_bbLoadOffsets_10 : _GEN_179; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_181 = 4'hb == _T_2014 ? io_bbLoadOffsets_11 : _GEN_180; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_182 = 4'hc == _T_2014 ? io_bbLoadOffsets_12 : _GEN_181; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_183 = 4'hd == _T_2014 ? io_bbLoadOffsets_13 : _GEN_182; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_184 = 4'he == _T_2014 ? io_bbLoadOffsets_14 : _GEN_183; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_185 = 4'hf == _T_2014 ? io_bbLoadOffsets_15 : _GEN_184; // @[LoadQueue.scala 77:20:@7934.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[LoadQueue.scala 76:25:@7927.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[LoadQueue.scala 76:25:@7927.4]
  assign _T_2032 = _T_1773[3:0]; // @[:@7949.6]
  assign _GEN_205 = 4'h1 == _T_2032 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_206 = 4'h2 == _T_2032 ? io_bbLoadOffsets_2 : _GEN_205; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_207 = 4'h3 == _T_2032 ? io_bbLoadOffsets_3 : _GEN_206; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_208 = 4'h4 == _T_2032 ? io_bbLoadOffsets_4 : _GEN_207; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_209 = 4'h5 == _T_2032 ? io_bbLoadOffsets_5 : _GEN_208; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_210 = 4'h6 == _T_2032 ? io_bbLoadOffsets_6 : _GEN_209; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_211 = 4'h7 == _T_2032 ? io_bbLoadOffsets_7 : _GEN_210; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_212 = 4'h8 == _T_2032 ? io_bbLoadOffsets_8 : _GEN_211; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_213 = 4'h9 == _T_2032 ? io_bbLoadOffsets_9 : _GEN_212; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_214 = 4'ha == _T_2032 ? io_bbLoadOffsets_10 : _GEN_213; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_215 = 4'hb == _T_2032 ? io_bbLoadOffsets_11 : _GEN_214; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_216 = 4'hc == _T_2032 ? io_bbLoadOffsets_12 : _GEN_215; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_217 = 4'hd == _T_2032 ? io_bbLoadOffsets_13 : _GEN_216; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_218 = 4'he == _T_2032 ? io_bbLoadOffsets_14 : _GEN_217; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_219 = 4'hf == _T_2032 ? io_bbLoadOffsets_15 : _GEN_218; // @[LoadQueue.scala 77:20:@7950.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[LoadQueue.scala 76:25:@7943.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[LoadQueue.scala 76:25:@7943.4]
  assign _T_2050 = _T_1782[3:0]; // @[:@7965.6]
  assign _GEN_239 = 4'h1 == _T_2050 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_240 = 4'h2 == _T_2050 ? io_bbLoadOffsets_2 : _GEN_239; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_241 = 4'h3 == _T_2050 ? io_bbLoadOffsets_3 : _GEN_240; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_242 = 4'h4 == _T_2050 ? io_bbLoadOffsets_4 : _GEN_241; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_243 = 4'h5 == _T_2050 ? io_bbLoadOffsets_5 : _GEN_242; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_244 = 4'h6 == _T_2050 ? io_bbLoadOffsets_6 : _GEN_243; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_245 = 4'h7 == _T_2050 ? io_bbLoadOffsets_7 : _GEN_244; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_246 = 4'h8 == _T_2050 ? io_bbLoadOffsets_8 : _GEN_245; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_247 = 4'h9 == _T_2050 ? io_bbLoadOffsets_9 : _GEN_246; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_248 = 4'ha == _T_2050 ? io_bbLoadOffsets_10 : _GEN_247; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_249 = 4'hb == _T_2050 ? io_bbLoadOffsets_11 : _GEN_248; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_250 = 4'hc == _T_2050 ? io_bbLoadOffsets_12 : _GEN_249; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_251 = 4'hd == _T_2050 ? io_bbLoadOffsets_13 : _GEN_250; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_252 = 4'he == _T_2050 ? io_bbLoadOffsets_14 : _GEN_251; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_253 = 4'hf == _T_2050 ? io_bbLoadOffsets_15 : _GEN_252; // @[LoadQueue.scala 77:20:@7966.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[LoadQueue.scala 76:25:@7959.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[LoadQueue.scala 76:25:@7959.4]
  assign _T_2068 = _T_1791[3:0]; // @[:@7981.6]
  assign _GEN_273 = 4'h1 == _T_2068 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_274 = 4'h2 == _T_2068 ? io_bbLoadOffsets_2 : _GEN_273; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_275 = 4'h3 == _T_2068 ? io_bbLoadOffsets_3 : _GEN_274; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_276 = 4'h4 == _T_2068 ? io_bbLoadOffsets_4 : _GEN_275; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_277 = 4'h5 == _T_2068 ? io_bbLoadOffsets_5 : _GEN_276; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_278 = 4'h6 == _T_2068 ? io_bbLoadOffsets_6 : _GEN_277; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_279 = 4'h7 == _T_2068 ? io_bbLoadOffsets_7 : _GEN_278; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_280 = 4'h8 == _T_2068 ? io_bbLoadOffsets_8 : _GEN_279; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_281 = 4'h9 == _T_2068 ? io_bbLoadOffsets_9 : _GEN_280; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_282 = 4'ha == _T_2068 ? io_bbLoadOffsets_10 : _GEN_281; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_283 = 4'hb == _T_2068 ? io_bbLoadOffsets_11 : _GEN_282; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_284 = 4'hc == _T_2068 ? io_bbLoadOffsets_12 : _GEN_283; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_285 = 4'hd == _T_2068 ? io_bbLoadOffsets_13 : _GEN_284; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_286 = 4'he == _T_2068 ? io_bbLoadOffsets_14 : _GEN_285; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_287 = 4'hf == _T_2068 ? io_bbLoadOffsets_15 : _GEN_286; // @[LoadQueue.scala 77:20:@7982.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[LoadQueue.scala 76:25:@7975.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[LoadQueue.scala 76:25:@7975.4]
  assign _T_2086 = _T_1800[3:0]; // @[:@7997.6]
  assign _GEN_307 = 4'h1 == _T_2086 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_308 = 4'h2 == _T_2086 ? io_bbLoadOffsets_2 : _GEN_307; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_309 = 4'h3 == _T_2086 ? io_bbLoadOffsets_3 : _GEN_308; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_310 = 4'h4 == _T_2086 ? io_bbLoadOffsets_4 : _GEN_309; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_311 = 4'h5 == _T_2086 ? io_bbLoadOffsets_5 : _GEN_310; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_312 = 4'h6 == _T_2086 ? io_bbLoadOffsets_6 : _GEN_311; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_313 = 4'h7 == _T_2086 ? io_bbLoadOffsets_7 : _GEN_312; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_314 = 4'h8 == _T_2086 ? io_bbLoadOffsets_8 : _GEN_313; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_315 = 4'h9 == _T_2086 ? io_bbLoadOffsets_9 : _GEN_314; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_316 = 4'ha == _T_2086 ? io_bbLoadOffsets_10 : _GEN_315; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_317 = 4'hb == _T_2086 ? io_bbLoadOffsets_11 : _GEN_316; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_318 = 4'hc == _T_2086 ? io_bbLoadOffsets_12 : _GEN_317; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_319 = 4'hd == _T_2086 ? io_bbLoadOffsets_13 : _GEN_318; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_320 = 4'he == _T_2086 ? io_bbLoadOffsets_14 : _GEN_319; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_321 = 4'hf == _T_2086 ? io_bbLoadOffsets_15 : _GEN_320; // @[LoadQueue.scala 77:20:@7998.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[LoadQueue.scala 76:25:@7991.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[LoadQueue.scala 76:25:@7991.4]
  assign _T_2104 = _T_1809[3:0]; // @[:@8013.6]
  assign _GEN_341 = 4'h1 == _T_2104 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_342 = 4'h2 == _T_2104 ? io_bbLoadOffsets_2 : _GEN_341; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_343 = 4'h3 == _T_2104 ? io_bbLoadOffsets_3 : _GEN_342; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_344 = 4'h4 == _T_2104 ? io_bbLoadOffsets_4 : _GEN_343; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_345 = 4'h5 == _T_2104 ? io_bbLoadOffsets_5 : _GEN_344; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_346 = 4'h6 == _T_2104 ? io_bbLoadOffsets_6 : _GEN_345; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_347 = 4'h7 == _T_2104 ? io_bbLoadOffsets_7 : _GEN_346; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_348 = 4'h8 == _T_2104 ? io_bbLoadOffsets_8 : _GEN_347; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_349 = 4'h9 == _T_2104 ? io_bbLoadOffsets_9 : _GEN_348; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_350 = 4'ha == _T_2104 ? io_bbLoadOffsets_10 : _GEN_349; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_351 = 4'hb == _T_2104 ? io_bbLoadOffsets_11 : _GEN_350; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_352 = 4'hc == _T_2104 ? io_bbLoadOffsets_12 : _GEN_351; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_353 = 4'hd == _T_2104 ? io_bbLoadOffsets_13 : _GEN_352; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_354 = 4'he == _T_2104 ? io_bbLoadOffsets_14 : _GEN_353; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_355 = 4'hf == _T_2104 ? io_bbLoadOffsets_15 : _GEN_354; // @[LoadQueue.scala 77:20:@8014.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[LoadQueue.scala 76:25:@8007.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[LoadQueue.scala 76:25:@8007.4]
  assign _T_2122 = _T_1818[3:0]; // @[:@8029.6]
  assign _GEN_375 = 4'h1 == _T_2122 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_376 = 4'h2 == _T_2122 ? io_bbLoadOffsets_2 : _GEN_375; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_377 = 4'h3 == _T_2122 ? io_bbLoadOffsets_3 : _GEN_376; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_378 = 4'h4 == _T_2122 ? io_bbLoadOffsets_4 : _GEN_377; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_379 = 4'h5 == _T_2122 ? io_bbLoadOffsets_5 : _GEN_378; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_380 = 4'h6 == _T_2122 ? io_bbLoadOffsets_6 : _GEN_379; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_381 = 4'h7 == _T_2122 ? io_bbLoadOffsets_7 : _GEN_380; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_382 = 4'h8 == _T_2122 ? io_bbLoadOffsets_8 : _GEN_381; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_383 = 4'h9 == _T_2122 ? io_bbLoadOffsets_9 : _GEN_382; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_384 = 4'ha == _T_2122 ? io_bbLoadOffsets_10 : _GEN_383; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_385 = 4'hb == _T_2122 ? io_bbLoadOffsets_11 : _GEN_384; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_386 = 4'hc == _T_2122 ? io_bbLoadOffsets_12 : _GEN_385; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_387 = 4'hd == _T_2122 ? io_bbLoadOffsets_13 : _GEN_386; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_388 = 4'he == _T_2122 ? io_bbLoadOffsets_14 : _GEN_387; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_389 = 4'hf == _T_2122 ? io_bbLoadOffsets_15 : _GEN_388; // @[LoadQueue.scala 77:20:@8030.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[LoadQueue.scala 76:25:@8023.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[LoadQueue.scala 76:25:@8023.4]
  assign _T_2140 = _T_1827[3:0]; // @[:@8045.6]
  assign _GEN_409 = 4'h1 == _T_2140 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_410 = 4'h2 == _T_2140 ? io_bbLoadOffsets_2 : _GEN_409; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_411 = 4'h3 == _T_2140 ? io_bbLoadOffsets_3 : _GEN_410; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_412 = 4'h4 == _T_2140 ? io_bbLoadOffsets_4 : _GEN_411; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_413 = 4'h5 == _T_2140 ? io_bbLoadOffsets_5 : _GEN_412; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_414 = 4'h6 == _T_2140 ? io_bbLoadOffsets_6 : _GEN_413; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_415 = 4'h7 == _T_2140 ? io_bbLoadOffsets_7 : _GEN_414; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_416 = 4'h8 == _T_2140 ? io_bbLoadOffsets_8 : _GEN_415; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_417 = 4'h9 == _T_2140 ? io_bbLoadOffsets_9 : _GEN_416; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_418 = 4'ha == _T_2140 ? io_bbLoadOffsets_10 : _GEN_417; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_419 = 4'hb == _T_2140 ? io_bbLoadOffsets_11 : _GEN_418; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_420 = 4'hc == _T_2140 ? io_bbLoadOffsets_12 : _GEN_419; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_421 = 4'hd == _T_2140 ? io_bbLoadOffsets_13 : _GEN_420; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_422 = 4'he == _T_2140 ? io_bbLoadOffsets_14 : _GEN_421; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_423 = 4'hf == _T_2140 ? io_bbLoadOffsets_15 : _GEN_422; // @[LoadQueue.scala 77:20:@8046.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[LoadQueue.scala 76:25:@8039.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[LoadQueue.scala 76:25:@8039.4]
  assign _T_2158 = _T_1836[3:0]; // @[:@8061.6]
  assign _GEN_443 = 4'h1 == _T_2158 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_444 = 4'h2 == _T_2158 ? io_bbLoadOffsets_2 : _GEN_443; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_445 = 4'h3 == _T_2158 ? io_bbLoadOffsets_3 : _GEN_444; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_446 = 4'h4 == _T_2158 ? io_bbLoadOffsets_4 : _GEN_445; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_447 = 4'h5 == _T_2158 ? io_bbLoadOffsets_5 : _GEN_446; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_448 = 4'h6 == _T_2158 ? io_bbLoadOffsets_6 : _GEN_447; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_449 = 4'h7 == _T_2158 ? io_bbLoadOffsets_7 : _GEN_448; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_450 = 4'h8 == _T_2158 ? io_bbLoadOffsets_8 : _GEN_449; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_451 = 4'h9 == _T_2158 ? io_bbLoadOffsets_9 : _GEN_450; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_452 = 4'ha == _T_2158 ? io_bbLoadOffsets_10 : _GEN_451; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_453 = 4'hb == _T_2158 ? io_bbLoadOffsets_11 : _GEN_452; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_454 = 4'hc == _T_2158 ? io_bbLoadOffsets_12 : _GEN_453; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_455 = 4'hd == _T_2158 ? io_bbLoadOffsets_13 : _GEN_454; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_456 = 4'he == _T_2158 ? io_bbLoadOffsets_14 : _GEN_455; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_457 = 4'hf == _T_2158 ? io_bbLoadOffsets_15 : _GEN_456; // @[LoadQueue.scala 77:20:@8062.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[LoadQueue.scala 76:25:@8055.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[LoadQueue.scala 76:25:@8055.4]
  assign _T_2176 = _T_1845[3:0]; // @[:@8077.6]
  assign _GEN_477 = 4'h1 == _T_2176 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_478 = 4'h2 == _T_2176 ? io_bbLoadOffsets_2 : _GEN_477; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_479 = 4'h3 == _T_2176 ? io_bbLoadOffsets_3 : _GEN_478; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_480 = 4'h4 == _T_2176 ? io_bbLoadOffsets_4 : _GEN_479; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_481 = 4'h5 == _T_2176 ? io_bbLoadOffsets_5 : _GEN_480; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_482 = 4'h6 == _T_2176 ? io_bbLoadOffsets_6 : _GEN_481; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_483 = 4'h7 == _T_2176 ? io_bbLoadOffsets_7 : _GEN_482; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_484 = 4'h8 == _T_2176 ? io_bbLoadOffsets_8 : _GEN_483; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_485 = 4'h9 == _T_2176 ? io_bbLoadOffsets_9 : _GEN_484; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_486 = 4'ha == _T_2176 ? io_bbLoadOffsets_10 : _GEN_485; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_487 = 4'hb == _T_2176 ? io_bbLoadOffsets_11 : _GEN_486; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_488 = 4'hc == _T_2176 ? io_bbLoadOffsets_12 : _GEN_487; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_489 = 4'hd == _T_2176 ? io_bbLoadOffsets_13 : _GEN_488; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_490 = 4'he == _T_2176 ? io_bbLoadOffsets_14 : _GEN_489; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_491 = 4'hf == _T_2176 ? io_bbLoadOffsets_15 : _GEN_490; // @[LoadQueue.scala 77:20:@8078.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[LoadQueue.scala 76:25:@8071.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[LoadQueue.scala 76:25:@8071.4]
  assign _T_2194 = _T_1854[3:0]; // @[:@8093.6]
  assign _GEN_511 = 4'h1 == _T_2194 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_512 = 4'h2 == _T_2194 ? io_bbLoadOffsets_2 : _GEN_511; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_513 = 4'h3 == _T_2194 ? io_bbLoadOffsets_3 : _GEN_512; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_514 = 4'h4 == _T_2194 ? io_bbLoadOffsets_4 : _GEN_513; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_515 = 4'h5 == _T_2194 ? io_bbLoadOffsets_5 : _GEN_514; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_516 = 4'h6 == _T_2194 ? io_bbLoadOffsets_6 : _GEN_515; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_517 = 4'h7 == _T_2194 ? io_bbLoadOffsets_7 : _GEN_516; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_518 = 4'h8 == _T_2194 ? io_bbLoadOffsets_8 : _GEN_517; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_519 = 4'h9 == _T_2194 ? io_bbLoadOffsets_9 : _GEN_518; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_520 = 4'ha == _T_2194 ? io_bbLoadOffsets_10 : _GEN_519; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_521 = 4'hb == _T_2194 ? io_bbLoadOffsets_11 : _GEN_520; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_522 = 4'hc == _T_2194 ? io_bbLoadOffsets_12 : _GEN_521; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_523 = 4'hd == _T_2194 ? io_bbLoadOffsets_13 : _GEN_522; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_524 = 4'he == _T_2194 ? io_bbLoadOffsets_14 : _GEN_523; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_525 = 4'hf == _T_2194 ? io_bbLoadOffsets_15 : _GEN_524; // @[LoadQueue.scala 77:20:@8094.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[LoadQueue.scala 76:25:@8087.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[LoadQueue.scala 76:25:@8087.4]
  assign _T_2216 = _GEN_15 + 4'h1; // @[util.scala 10:8:@8112.6]
  assign _GEN_31 = _T_2216 % 5'h10; // @[util.scala 10:14:@8113.6]
  assign _T_2217 = _GEN_31[4:0]; // @[util.scala 10:14:@8113.6]
  assign _GEN_2327 = {{1'd0}, io_storeTail}; // @[LoadQueue.scala 97:56:@8114.6]
  assign _T_2218 = _T_2217 == _GEN_2327; // @[LoadQueue.scala 97:56:@8114.6]
  assign _T_2219 = io_storeEmpty & _T_2218; // @[LoadQueue.scala 96:50:@8115.6]
  assign _T_2221 = _T_2219 == 1'h0; // @[LoadQueue.scala 96:34:@8116.6]
  assign _T_2223 = previousStoreHead <= offsetQ_0; // @[LoadQueue.scala 101:36:@8124.8]
  assign _T_2224 = offsetQ_0 < io_storeHead; // @[LoadQueue.scala 101:86:@8125.8]
  assign _T_2225 = _T_2223 & _T_2224; // @[LoadQueue.scala 101:61:@8126.8]
  assign _T_2227 = previousStoreHead > io_storeHead; // @[LoadQueue.scala 103:36:@8131.10]
  assign _T_2228 = io_storeHead <= offsetQ_0; // @[LoadQueue.scala 103:69:@8132.10]
  assign _T_2229 = offsetQ_0 < previousStoreHead; // @[LoadQueue.scala 104:31:@8133.10]
  assign _T_2230 = _T_2228 & _T_2229; // @[LoadQueue.scala 103:94:@8134.10]
  assign _T_2232 = _T_2230 == 1'h0; // @[LoadQueue.scala 103:54:@8135.10]
  assign _T_2233 = _T_2227 & _T_2232; // @[LoadQueue.scala 103:51:@8136.10]
  assign _GEN_560 = _T_2233 ? 1'h0 : checkBits_0; // @[LoadQueue.scala 104:53:@8137.10]
  assign _GEN_561 = _T_2225 ? 1'h0 : _GEN_560; // @[LoadQueue.scala 101:102:@8127.8]
  assign _GEN_562 = io_storeEmpty ? 1'h0 : _GEN_561; // @[LoadQueue.scala 99:27:@8120.6]
  assign _GEN_563 = initBits_0 ? _T_2221 : _GEN_562; // @[LoadQueue.scala 95:34:@8105.4]
  assign _T_2246 = _GEN_49 + 4'h1; // @[util.scala 10:8:@8148.6]
  assign _GEN_34 = _T_2246 % 5'h10; // @[util.scala 10:14:@8149.6]
  assign _T_2247 = _GEN_34[4:0]; // @[util.scala 10:14:@8149.6]
  assign _T_2248 = _T_2247 == _GEN_2327; // @[LoadQueue.scala 97:56:@8150.6]
  assign _T_2249 = io_storeEmpty & _T_2248; // @[LoadQueue.scala 96:50:@8151.6]
  assign _T_2251 = _T_2249 == 1'h0; // @[LoadQueue.scala 96:34:@8152.6]
  assign _T_2253 = previousStoreHead <= offsetQ_1; // @[LoadQueue.scala 101:36:@8160.8]
  assign _T_2254 = offsetQ_1 < io_storeHead; // @[LoadQueue.scala 101:86:@8161.8]
  assign _T_2255 = _T_2253 & _T_2254; // @[LoadQueue.scala 101:61:@8162.8]
  assign _T_2258 = io_storeHead <= offsetQ_1; // @[LoadQueue.scala 103:69:@8168.10]
  assign _T_2259 = offsetQ_1 < previousStoreHead; // @[LoadQueue.scala 104:31:@8169.10]
  assign _T_2260 = _T_2258 & _T_2259; // @[LoadQueue.scala 103:94:@8170.10]
  assign _T_2262 = _T_2260 == 1'h0; // @[LoadQueue.scala 103:54:@8171.10]
  assign _T_2263 = _T_2227 & _T_2262; // @[LoadQueue.scala 103:51:@8172.10]
  assign _GEN_580 = _T_2263 ? 1'h0 : checkBits_1; // @[LoadQueue.scala 104:53:@8173.10]
  assign _GEN_581 = _T_2255 ? 1'h0 : _GEN_580; // @[LoadQueue.scala 101:102:@8163.8]
  assign _GEN_582 = io_storeEmpty ? 1'h0 : _GEN_581; // @[LoadQueue.scala 99:27:@8156.6]
  assign _GEN_583 = initBits_1 ? _T_2251 : _GEN_582; // @[LoadQueue.scala 95:34:@8141.4]
  assign _T_2276 = _GEN_83 + 4'h1; // @[util.scala 10:8:@8184.6]
  assign _GEN_50 = _T_2276 % 5'h10; // @[util.scala 10:14:@8185.6]
  assign _T_2277 = _GEN_50[4:0]; // @[util.scala 10:14:@8185.6]
  assign _T_2278 = _T_2277 == _GEN_2327; // @[LoadQueue.scala 97:56:@8186.6]
  assign _T_2279 = io_storeEmpty & _T_2278; // @[LoadQueue.scala 96:50:@8187.6]
  assign _T_2281 = _T_2279 == 1'h0; // @[LoadQueue.scala 96:34:@8188.6]
  assign _T_2283 = previousStoreHead <= offsetQ_2; // @[LoadQueue.scala 101:36:@8196.8]
  assign _T_2284 = offsetQ_2 < io_storeHead; // @[LoadQueue.scala 101:86:@8197.8]
  assign _T_2285 = _T_2283 & _T_2284; // @[LoadQueue.scala 101:61:@8198.8]
  assign _T_2288 = io_storeHead <= offsetQ_2; // @[LoadQueue.scala 103:69:@8204.10]
  assign _T_2289 = offsetQ_2 < previousStoreHead; // @[LoadQueue.scala 104:31:@8205.10]
  assign _T_2290 = _T_2288 & _T_2289; // @[LoadQueue.scala 103:94:@8206.10]
  assign _T_2292 = _T_2290 == 1'h0; // @[LoadQueue.scala 103:54:@8207.10]
  assign _T_2293 = _T_2227 & _T_2292; // @[LoadQueue.scala 103:51:@8208.10]
  assign _GEN_600 = _T_2293 ? 1'h0 : checkBits_2; // @[LoadQueue.scala 104:53:@8209.10]
  assign _GEN_601 = _T_2285 ? 1'h0 : _GEN_600; // @[LoadQueue.scala 101:102:@8199.8]
  assign _GEN_602 = io_storeEmpty ? 1'h0 : _GEN_601; // @[LoadQueue.scala 99:27:@8192.6]
  assign _GEN_603 = initBits_2 ? _T_2281 : _GEN_602; // @[LoadQueue.scala 95:34:@8177.4]
  assign _T_2306 = _GEN_117 + 4'h1; // @[util.scala 10:8:@8220.6]
  assign _GEN_51 = _T_2306 % 5'h10; // @[util.scala 10:14:@8221.6]
  assign _T_2307 = _GEN_51[4:0]; // @[util.scala 10:14:@8221.6]
  assign _T_2308 = _T_2307 == _GEN_2327; // @[LoadQueue.scala 97:56:@8222.6]
  assign _T_2309 = io_storeEmpty & _T_2308; // @[LoadQueue.scala 96:50:@8223.6]
  assign _T_2311 = _T_2309 == 1'h0; // @[LoadQueue.scala 96:34:@8224.6]
  assign _T_2313 = previousStoreHead <= offsetQ_3; // @[LoadQueue.scala 101:36:@8232.8]
  assign _T_2314 = offsetQ_3 < io_storeHead; // @[LoadQueue.scala 101:86:@8233.8]
  assign _T_2315 = _T_2313 & _T_2314; // @[LoadQueue.scala 101:61:@8234.8]
  assign _T_2318 = io_storeHead <= offsetQ_3; // @[LoadQueue.scala 103:69:@8240.10]
  assign _T_2319 = offsetQ_3 < previousStoreHead; // @[LoadQueue.scala 104:31:@8241.10]
  assign _T_2320 = _T_2318 & _T_2319; // @[LoadQueue.scala 103:94:@8242.10]
  assign _T_2322 = _T_2320 == 1'h0; // @[LoadQueue.scala 103:54:@8243.10]
  assign _T_2323 = _T_2227 & _T_2322; // @[LoadQueue.scala 103:51:@8244.10]
  assign _GEN_620 = _T_2323 ? 1'h0 : checkBits_3; // @[LoadQueue.scala 104:53:@8245.10]
  assign _GEN_621 = _T_2315 ? 1'h0 : _GEN_620; // @[LoadQueue.scala 101:102:@8235.8]
  assign _GEN_622 = io_storeEmpty ? 1'h0 : _GEN_621; // @[LoadQueue.scala 99:27:@8228.6]
  assign _GEN_623 = initBits_3 ? _T_2311 : _GEN_622; // @[LoadQueue.scala 95:34:@8213.4]
  assign _T_2336 = _GEN_151 + 4'h1; // @[util.scala 10:8:@8256.6]
  assign _GEN_52 = _T_2336 % 5'h10; // @[util.scala 10:14:@8257.6]
  assign _T_2337 = _GEN_52[4:0]; // @[util.scala 10:14:@8257.6]
  assign _T_2338 = _T_2337 == _GEN_2327; // @[LoadQueue.scala 97:56:@8258.6]
  assign _T_2339 = io_storeEmpty & _T_2338; // @[LoadQueue.scala 96:50:@8259.6]
  assign _T_2341 = _T_2339 == 1'h0; // @[LoadQueue.scala 96:34:@8260.6]
  assign _T_2343 = previousStoreHead <= offsetQ_4; // @[LoadQueue.scala 101:36:@8268.8]
  assign _T_2344 = offsetQ_4 < io_storeHead; // @[LoadQueue.scala 101:86:@8269.8]
  assign _T_2345 = _T_2343 & _T_2344; // @[LoadQueue.scala 101:61:@8270.8]
  assign _T_2348 = io_storeHead <= offsetQ_4; // @[LoadQueue.scala 103:69:@8276.10]
  assign _T_2349 = offsetQ_4 < previousStoreHead; // @[LoadQueue.scala 104:31:@8277.10]
  assign _T_2350 = _T_2348 & _T_2349; // @[LoadQueue.scala 103:94:@8278.10]
  assign _T_2352 = _T_2350 == 1'h0; // @[LoadQueue.scala 103:54:@8279.10]
  assign _T_2353 = _T_2227 & _T_2352; // @[LoadQueue.scala 103:51:@8280.10]
  assign _GEN_640 = _T_2353 ? 1'h0 : checkBits_4; // @[LoadQueue.scala 104:53:@8281.10]
  assign _GEN_641 = _T_2345 ? 1'h0 : _GEN_640; // @[LoadQueue.scala 101:102:@8271.8]
  assign _GEN_642 = io_storeEmpty ? 1'h0 : _GEN_641; // @[LoadQueue.scala 99:27:@8264.6]
  assign _GEN_643 = initBits_4 ? _T_2341 : _GEN_642; // @[LoadQueue.scala 95:34:@8249.4]
  assign _T_2366 = _GEN_185 + 4'h1; // @[util.scala 10:8:@8292.6]
  assign _GEN_53 = _T_2366 % 5'h10; // @[util.scala 10:14:@8293.6]
  assign _T_2367 = _GEN_53[4:0]; // @[util.scala 10:14:@8293.6]
  assign _T_2368 = _T_2367 == _GEN_2327; // @[LoadQueue.scala 97:56:@8294.6]
  assign _T_2369 = io_storeEmpty & _T_2368; // @[LoadQueue.scala 96:50:@8295.6]
  assign _T_2371 = _T_2369 == 1'h0; // @[LoadQueue.scala 96:34:@8296.6]
  assign _T_2373 = previousStoreHead <= offsetQ_5; // @[LoadQueue.scala 101:36:@8304.8]
  assign _T_2374 = offsetQ_5 < io_storeHead; // @[LoadQueue.scala 101:86:@8305.8]
  assign _T_2375 = _T_2373 & _T_2374; // @[LoadQueue.scala 101:61:@8306.8]
  assign _T_2378 = io_storeHead <= offsetQ_5; // @[LoadQueue.scala 103:69:@8312.10]
  assign _T_2379 = offsetQ_5 < previousStoreHead; // @[LoadQueue.scala 104:31:@8313.10]
  assign _T_2380 = _T_2378 & _T_2379; // @[LoadQueue.scala 103:94:@8314.10]
  assign _T_2382 = _T_2380 == 1'h0; // @[LoadQueue.scala 103:54:@8315.10]
  assign _T_2383 = _T_2227 & _T_2382; // @[LoadQueue.scala 103:51:@8316.10]
  assign _GEN_660 = _T_2383 ? 1'h0 : checkBits_5; // @[LoadQueue.scala 104:53:@8317.10]
  assign _GEN_661 = _T_2375 ? 1'h0 : _GEN_660; // @[LoadQueue.scala 101:102:@8307.8]
  assign _GEN_662 = io_storeEmpty ? 1'h0 : _GEN_661; // @[LoadQueue.scala 99:27:@8300.6]
  assign _GEN_663 = initBits_5 ? _T_2371 : _GEN_662; // @[LoadQueue.scala 95:34:@8285.4]
  assign _T_2396 = _GEN_219 + 4'h1; // @[util.scala 10:8:@8328.6]
  assign _GEN_54 = _T_2396 % 5'h10; // @[util.scala 10:14:@8329.6]
  assign _T_2397 = _GEN_54[4:0]; // @[util.scala 10:14:@8329.6]
  assign _T_2398 = _T_2397 == _GEN_2327; // @[LoadQueue.scala 97:56:@8330.6]
  assign _T_2399 = io_storeEmpty & _T_2398; // @[LoadQueue.scala 96:50:@8331.6]
  assign _T_2401 = _T_2399 == 1'h0; // @[LoadQueue.scala 96:34:@8332.6]
  assign _T_2403 = previousStoreHead <= offsetQ_6; // @[LoadQueue.scala 101:36:@8340.8]
  assign _T_2404 = offsetQ_6 < io_storeHead; // @[LoadQueue.scala 101:86:@8341.8]
  assign _T_2405 = _T_2403 & _T_2404; // @[LoadQueue.scala 101:61:@8342.8]
  assign _T_2408 = io_storeHead <= offsetQ_6; // @[LoadQueue.scala 103:69:@8348.10]
  assign _T_2409 = offsetQ_6 < previousStoreHead; // @[LoadQueue.scala 104:31:@8349.10]
  assign _T_2410 = _T_2408 & _T_2409; // @[LoadQueue.scala 103:94:@8350.10]
  assign _T_2412 = _T_2410 == 1'h0; // @[LoadQueue.scala 103:54:@8351.10]
  assign _T_2413 = _T_2227 & _T_2412; // @[LoadQueue.scala 103:51:@8352.10]
  assign _GEN_680 = _T_2413 ? 1'h0 : checkBits_6; // @[LoadQueue.scala 104:53:@8353.10]
  assign _GEN_681 = _T_2405 ? 1'h0 : _GEN_680; // @[LoadQueue.scala 101:102:@8343.8]
  assign _GEN_682 = io_storeEmpty ? 1'h0 : _GEN_681; // @[LoadQueue.scala 99:27:@8336.6]
  assign _GEN_683 = initBits_6 ? _T_2401 : _GEN_682; // @[LoadQueue.scala 95:34:@8321.4]
  assign _T_2426 = _GEN_253 + 4'h1; // @[util.scala 10:8:@8364.6]
  assign _GEN_55 = _T_2426 % 5'h10; // @[util.scala 10:14:@8365.6]
  assign _T_2427 = _GEN_55[4:0]; // @[util.scala 10:14:@8365.6]
  assign _T_2428 = _T_2427 == _GEN_2327; // @[LoadQueue.scala 97:56:@8366.6]
  assign _T_2429 = io_storeEmpty & _T_2428; // @[LoadQueue.scala 96:50:@8367.6]
  assign _T_2431 = _T_2429 == 1'h0; // @[LoadQueue.scala 96:34:@8368.6]
  assign _T_2433 = previousStoreHead <= offsetQ_7; // @[LoadQueue.scala 101:36:@8376.8]
  assign _T_2434 = offsetQ_7 < io_storeHead; // @[LoadQueue.scala 101:86:@8377.8]
  assign _T_2435 = _T_2433 & _T_2434; // @[LoadQueue.scala 101:61:@8378.8]
  assign _T_2438 = io_storeHead <= offsetQ_7; // @[LoadQueue.scala 103:69:@8384.10]
  assign _T_2439 = offsetQ_7 < previousStoreHead; // @[LoadQueue.scala 104:31:@8385.10]
  assign _T_2440 = _T_2438 & _T_2439; // @[LoadQueue.scala 103:94:@8386.10]
  assign _T_2442 = _T_2440 == 1'h0; // @[LoadQueue.scala 103:54:@8387.10]
  assign _T_2443 = _T_2227 & _T_2442; // @[LoadQueue.scala 103:51:@8388.10]
  assign _GEN_700 = _T_2443 ? 1'h0 : checkBits_7; // @[LoadQueue.scala 104:53:@8389.10]
  assign _GEN_701 = _T_2435 ? 1'h0 : _GEN_700; // @[LoadQueue.scala 101:102:@8379.8]
  assign _GEN_702 = io_storeEmpty ? 1'h0 : _GEN_701; // @[LoadQueue.scala 99:27:@8372.6]
  assign _GEN_703 = initBits_7 ? _T_2431 : _GEN_702; // @[LoadQueue.scala 95:34:@8357.4]
  assign _T_2456 = _GEN_287 + 4'h1; // @[util.scala 10:8:@8400.6]
  assign _GEN_56 = _T_2456 % 5'h10; // @[util.scala 10:14:@8401.6]
  assign _T_2457 = _GEN_56[4:0]; // @[util.scala 10:14:@8401.6]
  assign _T_2458 = _T_2457 == _GEN_2327; // @[LoadQueue.scala 97:56:@8402.6]
  assign _T_2459 = io_storeEmpty & _T_2458; // @[LoadQueue.scala 96:50:@8403.6]
  assign _T_2461 = _T_2459 == 1'h0; // @[LoadQueue.scala 96:34:@8404.6]
  assign _T_2463 = previousStoreHead <= offsetQ_8; // @[LoadQueue.scala 101:36:@8412.8]
  assign _T_2464 = offsetQ_8 < io_storeHead; // @[LoadQueue.scala 101:86:@8413.8]
  assign _T_2465 = _T_2463 & _T_2464; // @[LoadQueue.scala 101:61:@8414.8]
  assign _T_2468 = io_storeHead <= offsetQ_8; // @[LoadQueue.scala 103:69:@8420.10]
  assign _T_2469 = offsetQ_8 < previousStoreHead; // @[LoadQueue.scala 104:31:@8421.10]
  assign _T_2470 = _T_2468 & _T_2469; // @[LoadQueue.scala 103:94:@8422.10]
  assign _T_2472 = _T_2470 == 1'h0; // @[LoadQueue.scala 103:54:@8423.10]
  assign _T_2473 = _T_2227 & _T_2472; // @[LoadQueue.scala 103:51:@8424.10]
  assign _GEN_720 = _T_2473 ? 1'h0 : checkBits_8; // @[LoadQueue.scala 104:53:@8425.10]
  assign _GEN_721 = _T_2465 ? 1'h0 : _GEN_720; // @[LoadQueue.scala 101:102:@8415.8]
  assign _GEN_722 = io_storeEmpty ? 1'h0 : _GEN_721; // @[LoadQueue.scala 99:27:@8408.6]
  assign _GEN_723 = initBits_8 ? _T_2461 : _GEN_722; // @[LoadQueue.scala 95:34:@8393.4]
  assign _T_2486 = _GEN_321 + 4'h1; // @[util.scala 10:8:@8436.6]
  assign _GEN_57 = _T_2486 % 5'h10; // @[util.scala 10:14:@8437.6]
  assign _T_2487 = _GEN_57[4:0]; // @[util.scala 10:14:@8437.6]
  assign _T_2488 = _T_2487 == _GEN_2327; // @[LoadQueue.scala 97:56:@8438.6]
  assign _T_2489 = io_storeEmpty & _T_2488; // @[LoadQueue.scala 96:50:@8439.6]
  assign _T_2491 = _T_2489 == 1'h0; // @[LoadQueue.scala 96:34:@8440.6]
  assign _T_2493 = previousStoreHead <= offsetQ_9; // @[LoadQueue.scala 101:36:@8448.8]
  assign _T_2494 = offsetQ_9 < io_storeHead; // @[LoadQueue.scala 101:86:@8449.8]
  assign _T_2495 = _T_2493 & _T_2494; // @[LoadQueue.scala 101:61:@8450.8]
  assign _T_2498 = io_storeHead <= offsetQ_9; // @[LoadQueue.scala 103:69:@8456.10]
  assign _T_2499 = offsetQ_9 < previousStoreHead; // @[LoadQueue.scala 104:31:@8457.10]
  assign _T_2500 = _T_2498 & _T_2499; // @[LoadQueue.scala 103:94:@8458.10]
  assign _T_2502 = _T_2500 == 1'h0; // @[LoadQueue.scala 103:54:@8459.10]
  assign _T_2503 = _T_2227 & _T_2502; // @[LoadQueue.scala 103:51:@8460.10]
  assign _GEN_740 = _T_2503 ? 1'h0 : checkBits_9; // @[LoadQueue.scala 104:53:@8461.10]
  assign _GEN_741 = _T_2495 ? 1'h0 : _GEN_740; // @[LoadQueue.scala 101:102:@8451.8]
  assign _GEN_742 = io_storeEmpty ? 1'h0 : _GEN_741; // @[LoadQueue.scala 99:27:@8444.6]
  assign _GEN_743 = initBits_9 ? _T_2491 : _GEN_742; // @[LoadQueue.scala 95:34:@8429.4]
  assign _T_2516 = _GEN_355 + 4'h1; // @[util.scala 10:8:@8472.6]
  assign _GEN_58 = _T_2516 % 5'h10; // @[util.scala 10:14:@8473.6]
  assign _T_2517 = _GEN_58[4:0]; // @[util.scala 10:14:@8473.6]
  assign _T_2518 = _T_2517 == _GEN_2327; // @[LoadQueue.scala 97:56:@8474.6]
  assign _T_2519 = io_storeEmpty & _T_2518; // @[LoadQueue.scala 96:50:@8475.6]
  assign _T_2521 = _T_2519 == 1'h0; // @[LoadQueue.scala 96:34:@8476.6]
  assign _T_2523 = previousStoreHead <= offsetQ_10; // @[LoadQueue.scala 101:36:@8484.8]
  assign _T_2524 = offsetQ_10 < io_storeHead; // @[LoadQueue.scala 101:86:@8485.8]
  assign _T_2525 = _T_2523 & _T_2524; // @[LoadQueue.scala 101:61:@8486.8]
  assign _T_2528 = io_storeHead <= offsetQ_10; // @[LoadQueue.scala 103:69:@8492.10]
  assign _T_2529 = offsetQ_10 < previousStoreHead; // @[LoadQueue.scala 104:31:@8493.10]
  assign _T_2530 = _T_2528 & _T_2529; // @[LoadQueue.scala 103:94:@8494.10]
  assign _T_2532 = _T_2530 == 1'h0; // @[LoadQueue.scala 103:54:@8495.10]
  assign _T_2533 = _T_2227 & _T_2532; // @[LoadQueue.scala 103:51:@8496.10]
  assign _GEN_760 = _T_2533 ? 1'h0 : checkBits_10; // @[LoadQueue.scala 104:53:@8497.10]
  assign _GEN_761 = _T_2525 ? 1'h0 : _GEN_760; // @[LoadQueue.scala 101:102:@8487.8]
  assign _GEN_762 = io_storeEmpty ? 1'h0 : _GEN_761; // @[LoadQueue.scala 99:27:@8480.6]
  assign _GEN_763 = initBits_10 ? _T_2521 : _GEN_762; // @[LoadQueue.scala 95:34:@8465.4]
  assign _T_2546 = _GEN_389 + 4'h1; // @[util.scala 10:8:@8508.6]
  assign _GEN_59 = _T_2546 % 5'h10; // @[util.scala 10:14:@8509.6]
  assign _T_2547 = _GEN_59[4:0]; // @[util.scala 10:14:@8509.6]
  assign _T_2548 = _T_2547 == _GEN_2327; // @[LoadQueue.scala 97:56:@8510.6]
  assign _T_2549 = io_storeEmpty & _T_2548; // @[LoadQueue.scala 96:50:@8511.6]
  assign _T_2551 = _T_2549 == 1'h0; // @[LoadQueue.scala 96:34:@8512.6]
  assign _T_2553 = previousStoreHead <= offsetQ_11; // @[LoadQueue.scala 101:36:@8520.8]
  assign _T_2554 = offsetQ_11 < io_storeHead; // @[LoadQueue.scala 101:86:@8521.8]
  assign _T_2555 = _T_2553 & _T_2554; // @[LoadQueue.scala 101:61:@8522.8]
  assign _T_2558 = io_storeHead <= offsetQ_11; // @[LoadQueue.scala 103:69:@8528.10]
  assign _T_2559 = offsetQ_11 < previousStoreHead; // @[LoadQueue.scala 104:31:@8529.10]
  assign _T_2560 = _T_2558 & _T_2559; // @[LoadQueue.scala 103:94:@8530.10]
  assign _T_2562 = _T_2560 == 1'h0; // @[LoadQueue.scala 103:54:@8531.10]
  assign _T_2563 = _T_2227 & _T_2562; // @[LoadQueue.scala 103:51:@8532.10]
  assign _GEN_780 = _T_2563 ? 1'h0 : checkBits_11; // @[LoadQueue.scala 104:53:@8533.10]
  assign _GEN_781 = _T_2555 ? 1'h0 : _GEN_780; // @[LoadQueue.scala 101:102:@8523.8]
  assign _GEN_782 = io_storeEmpty ? 1'h0 : _GEN_781; // @[LoadQueue.scala 99:27:@8516.6]
  assign _GEN_783 = initBits_11 ? _T_2551 : _GEN_782; // @[LoadQueue.scala 95:34:@8501.4]
  assign _T_2576 = _GEN_423 + 4'h1; // @[util.scala 10:8:@8544.6]
  assign _GEN_60 = _T_2576 % 5'h10; // @[util.scala 10:14:@8545.6]
  assign _T_2577 = _GEN_60[4:0]; // @[util.scala 10:14:@8545.6]
  assign _T_2578 = _T_2577 == _GEN_2327; // @[LoadQueue.scala 97:56:@8546.6]
  assign _T_2579 = io_storeEmpty & _T_2578; // @[LoadQueue.scala 96:50:@8547.6]
  assign _T_2581 = _T_2579 == 1'h0; // @[LoadQueue.scala 96:34:@8548.6]
  assign _T_2583 = previousStoreHead <= offsetQ_12; // @[LoadQueue.scala 101:36:@8556.8]
  assign _T_2584 = offsetQ_12 < io_storeHead; // @[LoadQueue.scala 101:86:@8557.8]
  assign _T_2585 = _T_2583 & _T_2584; // @[LoadQueue.scala 101:61:@8558.8]
  assign _T_2588 = io_storeHead <= offsetQ_12; // @[LoadQueue.scala 103:69:@8564.10]
  assign _T_2589 = offsetQ_12 < previousStoreHead; // @[LoadQueue.scala 104:31:@8565.10]
  assign _T_2590 = _T_2588 & _T_2589; // @[LoadQueue.scala 103:94:@8566.10]
  assign _T_2592 = _T_2590 == 1'h0; // @[LoadQueue.scala 103:54:@8567.10]
  assign _T_2593 = _T_2227 & _T_2592; // @[LoadQueue.scala 103:51:@8568.10]
  assign _GEN_800 = _T_2593 ? 1'h0 : checkBits_12; // @[LoadQueue.scala 104:53:@8569.10]
  assign _GEN_801 = _T_2585 ? 1'h0 : _GEN_800; // @[LoadQueue.scala 101:102:@8559.8]
  assign _GEN_802 = io_storeEmpty ? 1'h0 : _GEN_801; // @[LoadQueue.scala 99:27:@8552.6]
  assign _GEN_803 = initBits_12 ? _T_2581 : _GEN_802; // @[LoadQueue.scala 95:34:@8537.4]
  assign _T_2606 = _GEN_457 + 4'h1; // @[util.scala 10:8:@8580.6]
  assign _GEN_61 = _T_2606 % 5'h10; // @[util.scala 10:14:@8581.6]
  assign _T_2607 = _GEN_61[4:0]; // @[util.scala 10:14:@8581.6]
  assign _T_2608 = _T_2607 == _GEN_2327; // @[LoadQueue.scala 97:56:@8582.6]
  assign _T_2609 = io_storeEmpty & _T_2608; // @[LoadQueue.scala 96:50:@8583.6]
  assign _T_2611 = _T_2609 == 1'h0; // @[LoadQueue.scala 96:34:@8584.6]
  assign _T_2613 = previousStoreHead <= offsetQ_13; // @[LoadQueue.scala 101:36:@8592.8]
  assign _T_2614 = offsetQ_13 < io_storeHead; // @[LoadQueue.scala 101:86:@8593.8]
  assign _T_2615 = _T_2613 & _T_2614; // @[LoadQueue.scala 101:61:@8594.8]
  assign _T_2618 = io_storeHead <= offsetQ_13; // @[LoadQueue.scala 103:69:@8600.10]
  assign _T_2619 = offsetQ_13 < previousStoreHead; // @[LoadQueue.scala 104:31:@8601.10]
  assign _T_2620 = _T_2618 & _T_2619; // @[LoadQueue.scala 103:94:@8602.10]
  assign _T_2622 = _T_2620 == 1'h0; // @[LoadQueue.scala 103:54:@8603.10]
  assign _T_2623 = _T_2227 & _T_2622; // @[LoadQueue.scala 103:51:@8604.10]
  assign _GEN_820 = _T_2623 ? 1'h0 : checkBits_13; // @[LoadQueue.scala 104:53:@8605.10]
  assign _GEN_821 = _T_2615 ? 1'h0 : _GEN_820; // @[LoadQueue.scala 101:102:@8595.8]
  assign _GEN_822 = io_storeEmpty ? 1'h0 : _GEN_821; // @[LoadQueue.scala 99:27:@8588.6]
  assign _GEN_823 = initBits_13 ? _T_2611 : _GEN_822; // @[LoadQueue.scala 95:34:@8573.4]
  assign _T_2636 = _GEN_491 + 4'h1; // @[util.scala 10:8:@8616.6]
  assign _GEN_62 = _T_2636 % 5'h10; // @[util.scala 10:14:@8617.6]
  assign _T_2637 = _GEN_62[4:0]; // @[util.scala 10:14:@8617.6]
  assign _T_2638 = _T_2637 == _GEN_2327; // @[LoadQueue.scala 97:56:@8618.6]
  assign _T_2639 = io_storeEmpty & _T_2638; // @[LoadQueue.scala 96:50:@8619.6]
  assign _T_2641 = _T_2639 == 1'h0; // @[LoadQueue.scala 96:34:@8620.6]
  assign _T_2643 = previousStoreHead <= offsetQ_14; // @[LoadQueue.scala 101:36:@8628.8]
  assign _T_2644 = offsetQ_14 < io_storeHead; // @[LoadQueue.scala 101:86:@8629.8]
  assign _T_2645 = _T_2643 & _T_2644; // @[LoadQueue.scala 101:61:@8630.8]
  assign _T_2648 = io_storeHead <= offsetQ_14; // @[LoadQueue.scala 103:69:@8636.10]
  assign _T_2649 = offsetQ_14 < previousStoreHead; // @[LoadQueue.scala 104:31:@8637.10]
  assign _T_2650 = _T_2648 & _T_2649; // @[LoadQueue.scala 103:94:@8638.10]
  assign _T_2652 = _T_2650 == 1'h0; // @[LoadQueue.scala 103:54:@8639.10]
  assign _T_2653 = _T_2227 & _T_2652; // @[LoadQueue.scala 103:51:@8640.10]
  assign _GEN_840 = _T_2653 ? 1'h0 : checkBits_14; // @[LoadQueue.scala 104:53:@8641.10]
  assign _GEN_841 = _T_2645 ? 1'h0 : _GEN_840; // @[LoadQueue.scala 101:102:@8631.8]
  assign _GEN_842 = io_storeEmpty ? 1'h0 : _GEN_841; // @[LoadQueue.scala 99:27:@8624.6]
  assign _GEN_843 = initBits_14 ? _T_2641 : _GEN_842; // @[LoadQueue.scala 95:34:@8609.4]
  assign _T_2666 = _GEN_525 + 4'h1; // @[util.scala 10:8:@8652.6]
  assign _GEN_63 = _T_2666 % 5'h10; // @[util.scala 10:14:@8653.6]
  assign _T_2667 = _GEN_63[4:0]; // @[util.scala 10:14:@8653.6]
  assign _T_2668 = _T_2667 == _GEN_2327; // @[LoadQueue.scala 97:56:@8654.6]
  assign _T_2669 = io_storeEmpty & _T_2668; // @[LoadQueue.scala 96:50:@8655.6]
  assign _T_2671 = _T_2669 == 1'h0; // @[LoadQueue.scala 96:34:@8656.6]
  assign _T_2673 = previousStoreHead <= offsetQ_15; // @[LoadQueue.scala 101:36:@8664.8]
  assign _T_2674 = offsetQ_15 < io_storeHead; // @[LoadQueue.scala 101:86:@8665.8]
  assign _T_2675 = _T_2673 & _T_2674; // @[LoadQueue.scala 101:61:@8666.8]
  assign _T_2678 = io_storeHead <= offsetQ_15; // @[LoadQueue.scala 103:69:@8672.10]
  assign _T_2679 = offsetQ_15 < previousStoreHead; // @[LoadQueue.scala 104:31:@8673.10]
  assign _T_2680 = _T_2678 & _T_2679; // @[LoadQueue.scala 103:94:@8674.10]
  assign _T_2682 = _T_2680 == 1'h0; // @[LoadQueue.scala 103:54:@8675.10]
  assign _T_2683 = _T_2227 & _T_2682; // @[LoadQueue.scala 103:51:@8676.10]
  assign _GEN_860 = _T_2683 ? 1'h0 : checkBits_15; // @[LoadQueue.scala 104:53:@8677.10]
  assign _GEN_861 = _T_2675 ? 1'h0 : _GEN_860; // @[LoadQueue.scala 101:102:@8667.8]
  assign _GEN_862 = io_storeEmpty ? 1'h0 : _GEN_861; // @[LoadQueue.scala 99:27:@8660.6]
  assign _GEN_863 = initBits_15 ? _T_2671 : _GEN_862; // @[LoadQueue.scala 95:34:@8645.4]
  assign _T_2687 = 16'h1 << io_storeHead; // @[OneHot.scala 52:12:@8682.4]
  assign _T_2689 = _T_2687[0]; // @[util.scala 60:60:@8684.4]
  assign _T_2690 = _T_2687[1]; // @[util.scala 60:60:@8685.4]
  assign _T_2691 = _T_2687[2]; // @[util.scala 60:60:@8686.4]
  assign _T_2692 = _T_2687[3]; // @[util.scala 60:60:@8687.4]
  assign _T_2693 = _T_2687[4]; // @[util.scala 60:60:@8688.4]
  assign _T_2694 = _T_2687[5]; // @[util.scala 60:60:@8689.4]
  assign _T_2695 = _T_2687[6]; // @[util.scala 60:60:@8690.4]
  assign _T_2696 = _T_2687[7]; // @[util.scala 60:60:@8691.4]
  assign _T_2697 = _T_2687[8]; // @[util.scala 60:60:@8692.4]
  assign _T_2698 = _T_2687[9]; // @[util.scala 60:60:@8693.4]
  assign _T_2699 = _T_2687[10]; // @[util.scala 60:60:@8694.4]
  assign _T_2700 = _T_2687[11]; // @[util.scala 60:60:@8695.4]
  assign _T_2701 = _T_2687[12]; // @[util.scala 60:60:@8696.4]
  assign _T_2702 = _T_2687[13]; // @[util.scala 60:60:@8697.4]
  assign _T_2703 = _T_2687[14]; // @[util.scala 60:60:@8698.4]
  assign _T_2704 = _T_2687[15]; // @[util.scala 60:60:@8699.4]
  assign _T_4835 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@10223.4]
  assign _T_4842 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8}; // @[Mux.scala 19:72:@10230.4]
  assign _T_4843 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,_T_4835}; // @[Mux.scala 19:72:@10231.4]
  assign _T_4845 = _T_2689 ? _T_4843 : 512'h0; // @[Mux.scala 19:72:@10232.4]
  assign _T_4852 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@10239.4]
  assign _T_4859 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9}; // @[Mux.scala 19:72:@10246.4]
  assign _T_4860 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,_T_4852}; // @[Mux.scala 19:72:@10247.4]
  assign _T_4862 = _T_2690 ? _T_4860 : 512'h0; // @[Mux.scala 19:72:@10248.4]
  assign _T_4869 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@10255.4]
  assign _T_4876 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10}; // @[Mux.scala 19:72:@10262.4]
  assign _T_4877 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,_T_4869}; // @[Mux.scala 19:72:@10263.4]
  assign _T_4879 = _T_2691 ? _T_4877 : 512'h0; // @[Mux.scala 19:72:@10264.4]
  assign _T_4886 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@10271.4]
  assign _T_4893 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11}; // @[Mux.scala 19:72:@10278.4]
  assign _T_4894 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,_T_4886}; // @[Mux.scala 19:72:@10279.4]
  assign _T_4896 = _T_2692 ? _T_4894 : 512'h0; // @[Mux.scala 19:72:@10280.4]
  assign _T_4903 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@10287.4]
  assign _T_4910 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12}; // @[Mux.scala 19:72:@10294.4]
  assign _T_4911 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,_T_4903}; // @[Mux.scala 19:72:@10295.4]
  assign _T_4913 = _T_2693 ? _T_4911 : 512'h0; // @[Mux.scala 19:72:@10296.4]
  assign _T_4920 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@10303.4]
  assign _T_4927 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13}; // @[Mux.scala 19:72:@10310.4]
  assign _T_4928 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,_T_4920}; // @[Mux.scala 19:72:@10311.4]
  assign _T_4930 = _T_2694 ? _T_4928 : 512'h0; // @[Mux.scala 19:72:@10312.4]
  assign _T_4937 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@10319.4]
  assign _T_4944 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14}; // @[Mux.scala 19:72:@10326.4]
  assign _T_4945 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,_T_4937}; // @[Mux.scala 19:72:@10327.4]
  assign _T_4947 = _T_2695 ? _T_4945 : 512'h0; // @[Mux.scala 19:72:@10328.4]
  assign _T_4954 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7}; // @[Mux.scala 19:72:@10335.4]
  assign _T_4961 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15}; // @[Mux.scala 19:72:@10342.4]
  assign _T_4962 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,_T_4954}; // @[Mux.scala 19:72:@10343.4]
  assign _T_4964 = _T_2696 ? _T_4962 : 512'h0; // @[Mux.scala 19:72:@10344.4]
  assign _T_4979 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,_T_4842}; // @[Mux.scala 19:72:@10359.4]
  assign _T_4981 = _T_2697 ? _T_4979 : 512'h0; // @[Mux.scala 19:72:@10360.4]
  assign _T_4996 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,_T_4859}; // @[Mux.scala 19:72:@10375.4]
  assign _T_4998 = _T_2698 ? _T_4996 : 512'h0; // @[Mux.scala 19:72:@10376.4]
  assign _T_5013 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,_T_4876}; // @[Mux.scala 19:72:@10391.4]
  assign _T_5015 = _T_2699 ? _T_5013 : 512'h0; // @[Mux.scala 19:72:@10392.4]
  assign _T_5030 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,_T_4893}; // @[Mux.scala 19:72:@10407.4]
  assign _T_5032 = _T_2700 ? _T_5030 : 512'h0; // @[Mux.scala 19:72:@10408.4]
  assign _T_5047 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,_T_4910}; // @[Mux.scala 19:72:@10423.4]
  assign _T_5049 = _T_2701 ? _T_5047 : 512'h0; // @[Mux.scala 19:72:@10424.4]
  assign _T_5064 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,_T_4927}; // @[Mux.scala 19:72:@10439.4]
  assign _T_5066 = _T_2702 ? _T_5064 : 512'h0; // @[Mux.scala 19:72:@10440.4]
  assign _T_5081 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,_T_4944}; // @[Mux.scala 19:72:@10455.4]
  assign _T_5083 = _T_2703 ? _T_5081 : 512'h0; // @[Mux.scala 19:72:@10456.4]
  assign _T_5098 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,_T_4961}; // @[Mux.scala 19:72:@10471.4]
  assign _T_5100 = _T_2704 ? _T_5098 : 512'h0; // @[Mux.scala 19:72:@10472.4]
  assign _T_5101 = _T_4845 | _T_4862; // @[Mux.scala 19:72:@10473.4]
  assign _T_5102 = _T_5101 | _T_4879; // @[Mux.scala 19:72:@10474.4]
  assign _T_5103 = _T_5102 | _T_4896; // @[Mux.scala 19:72:@10475.4]
  assign _T_5104 = _T_5103 | _T_4913; // @[Mux.scala 19:72:@10476.4]
  assign _T_5105 = _T_5104 | _T_4930; // @[Mux.scala 19:72:@10477.4]
  assign _T_5106 = _T_5105 | _T_4947; // @[Mux.scala 19:72:@10478.4]
  assign _T_5107 = _T_5106 | _T_4964; // @[Mux.scala 19:72:@10479.4]
  assign _T_5108 = _T_5107 | _T_4981; // @[Mux.scala 19:72:@10480.4]
  assign _T_5109 = _T_5108 | _T_4998; // @[Mux.scala 19:72:@10481.4]
  assign _T_5110 = _T_5109 | _T_5015; // @[Mux.scala 19:72:@10482.4]
  assign _T_5111 = _T_5110 | _T_5032; // @[Mux.scala 19:72:@10483.4]
  assign _T_5112 = _T_5111 | _T_5049; // @[Mux.scala 19:72:@10484.4]
  assign _T_5113 = _T_5112 | _T_5066; // @[Mux.scala 19:72:@10485.4]
  assign _T_5114 = _T_5113 | _T_5083; // @[Mux.scala 19:72:@10486.4]
  assign _T_5115 = _T_5114 | _T_5100; // @[Mux.scala 19:72:@10487.4]
  assign _T_5692 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@10837.4]
  assign _T_5699 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8}; // @[Mux.scala 19:72:@10844.4]
  assign _T_5700 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,_T_5692}; // @[Mux.scala 19:72:@10845.4]
  assign _T_5702 = _T_2689 ? _T_5700 : 16'h0; // @[Mux.scala 19:72:@10846.4]
  assign _T_5709 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@10853.4]
  assign _T_5716 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9}; // @[Mux.scala 19:72:@10860.4]
  assign _T_5717 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,_T_5709}; // @[Mux.scala 19:72:@10861.4]
  assign _T_5719 = _T_2690 ? _T_5717 : 16'h0; // @[Mux.scala 19:72:@10862.4]
  assign _T_5726 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@10869.4]
  assign _T_5733 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10}; // @[Mux.scala 19:72:@10876.4]
  assign _T_5734 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,_T_5726}; // @[Mux.scala 19:72:@10877.4]
  assign _T_5736 = _T_2691 ? _T_5734 : 16'h0; // @[Mux.scala 19:72:@10878.4]
  assign _T_5743 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@10885.4]
  assign _T_5750 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11}; // @[Mux.scala 19:72:@10892.4]
  assign _T_5751 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,_T_5743}; // @[Mux.scala 19:72:@10893.4]
  assign _T_5753 = _T_2692 ? _T_5751 : 16'h0; // @[Mux.scala 19:72:@10894.4]
  assign _T_5760 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@10901.4]
  assign _T_5767 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12}; // @[Mux.scala 19:72:@10908.4]
  assign _T_5768 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,_T_5760}; // @[Mux.scala 19:72:@10909.4]
  assign _T_5770 = _T_2693 ? _T_5768 : 16'h0; // @[Mux.scala 19:72:@10910.4]
  assign _T_5777 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@10917.4]
  assign _T_5784 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13}; // @[Mux.scala 19:72:@10924.4]
  assign _T_5785 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,_T_5777}; // @[Mux.scala 19:72:@10925.4]
  assign _T_5787 = _T_2694 ? _T_5785 : 16'h0; // @[Mux.scala 19:72:@10926.4]
  assign _T_5794 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@10933.4]
  assign _T_5801 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14}; // @[Mux.scala 19:72:@10940.4]
  assign _T_5802 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,_T_5794}; // @[Mux.scala 19:72:@10941.4]
  assign _T_5804 = _T_2695 ? _T_5802 : 16'h0; // @[Mux.scala 19:72:@10942.4]
  assign _T_5811 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7}; // @[Mux.scala 19:72:@10949.4]
  assign _T_5818 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15}; // @[Mux.scala 19:72:@10956.4]
  assign _T_5819 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,_T_5811}; // @[Mux.scala 19:72:@10957.4]
  assign _T_5821 = _T_2696 ? _T_5819 : 16'h0; // @[Mux.scala 19:72:@10958.4]
  assign _T_5836 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,_T_5699}; // @[Mux.scala 19:72:@10973.4]
  assign _T_5838 = _T_2697 ? _T_5836 : 16'h0; // @[Mux.scala 19:72:@10974.4]
  assign _T_5853 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,_T_5716}; // @[Mux.scala 19:72:@10989.4]
  assign _T_5855 = _T_2698 ? _T_5853 : 16'h0; // @[Mux.scala 19:72:@10990.4]
  assign _T_5870 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,_T_5733}; // @[Mux.scala 19:72:@11005.4]
  assign _T_5872 = _T_2699 ? _T_5870 : 16'h0; // @[Mux.scala 19:72:@11006.4]
  assign _T_5887 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,_T_5750}; // @[Mux.scala 19:72:@11021.4]
  assign _T_5889 = _T_2700 ? _T_5887 : 16'h0; // @[Mux.scala 19:72:@11022.4]
  assign _T_5904 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,_T_5767}; // @[Mux.scala 19:72:@11037.4]
  assign _T_5906 = _T_2701 ? _T_5904 : 16'h0; // @[Mux.scala 19:72:@11038.4]
  assign _T_5921 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,_T_5784}; // @[Mux.scala 19:72:@11053.4]
  assign _T_5923 = _T_2702 ? _T_5921 : 16'h0; // @[Mux.scala 19:72:@11054.4]
  assign _T_5938 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,_T_5801}; // @[Mux.scala 19:72:@11069.4]
  assign _T_5940 = _T_2703 ? _T_5938 : 16'h0; // @[Mux.scala 19:72:@11070.4]
  assign _T_5955 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,_T_5818}; // @[Mux.scala 19:72:@11085.4]
  assign _T_5957 = _T_2704 ? _T_5955 : 16'h0; // @[Mux.scala 19:72:@11086.4]
  assign _T_5958 = _T_5702 | _T_5719; // @[Mux.scala 19:72:@11087.4]
  assign _T_5959 = _T_5958 | _T_5736; // @[Mux.scala 19:72:@11088.4]
  assign _T_5960 = _T_5959 | _T_5753; // @[Mux.scala 19:72:@11089.4]
  assign _T_5961 = _T_5960 | _T_5770; // @[Mux.scala 19:72:@11090.4]
  assign _T_5962 = _T_5961 | _T_5787; // @[Mux.scala 19:72:@11091.4]
  assign _T_5963 = _T_5962 | _T_5804; // @[Mux.scala 19:72:@11092.4]
  assign _T_5964 = _T_5963 | _T_5821; // @[Mux.scala 19:72:@11093.4]
  assign _T_5965 = _T_5964 | _T_5838; // @[Mux.scala 19:72:@11094.4]
  assign _T_5966 = _T_5965 | _T_5855; // @[Mux.scala 19:72:@11095.4]
  assign _T_5967 = _T_5966 | _T_5872; // @[Mux.scala 19:72:@11096.4]
  assign _T_5968 = _T_5967 | _T_5889; // @[Mux.scala 19:72:@11097.4]
  assign _T_5969 = _T_5968 | _T_5906; // @[Mux.scala 19:72:@11098.4]
  assign _T_5970 = _T_5969 | _T_5923; // @[Mux.scala 19:72:@11099.4]
  assign _T_5971 = _T_5970 | _T_5940; // @[Mux.scala 19:72:@11100.4]
  assign _T_5972 = _T_5971 | _T_5957; // @[Mux.scala 19:72:@11101.4]
  assign _T_6113 = io_storeHead < io_storeTail; // @[LoadQueue.scala 121:105:@11137.4]
  assign _T_6115 = io_storeHead <= 4'h0; // @[LoadQueue.scala 122:18:@11138.4]
  assign _T_6117 = 4'h0 < io_storeTail; // @[LoadQueue.scala 122:36:@11139.4]
  assign _T_6118 = _T_6115 & _T_6117; // @[LoadQueue.scala 122:27:@11140.4]
  assign _T_6120 = io_storeEmpty == 1'h0; // @[LoadQueue.scala 122:52:@11141.4]
  assign _T_6122 = io_storeTail <= 4'h0; // @[LoadQueue.scala 122:85:@11142.4]
  assign _T_6124 = 4'h0 < io_storeHead; // @[LoadQueue.scala 122:103:@11143.4]
  assign _T_6125 = _T_6122 & _T_6124; // @[LoadQueue.scala 122:94:@11144.4]
  assign _T_6127 = _T_6125 == 1'h0; // @[LoadQueue.scala 122:70:@11145.4]
  assign _T_6128 = _T_6120 & _T_6127; // @[LoadQueue.scala 122:67:@11146.4]
  assign validEntriesInStoreQ_0 = _T_6113 ? _T_6118 : _T_6128; // @[LoadQueue.scala 121:91:@11147.4]
  assign _T_6132 = io_storeHead <= 4'h1; // @[LoadQueue.scala 122:18:@11149.4]
  assign _T_6134 = 4'h1 < io_storeTail; // @[LoadQueue.scala 122:36:@11150.4]
  assign _T_6135 = _T_6132 & _T_6134; // @[LoadQueue.scala 122:27:@11151.4]
  assign _T_6139 = io_storeTail <= 4'h1; // @[LoadQueue.scala 122:85:@11153.4]
  assign _T_6141 = 4'h1 < io_storeHead; // @[LoadQueue.scala 122:103:@11154.4]
  assign _T_6142 = _T_6139 & _T_6141; // @[LoadQueue.scala 122:94:@11155.4]
  assign _T_6144 = _T_6142 == 1'h0; // @[LoadQueue.scala 122:70:@11156.4]
  assign _T_6145 = _T_6120 & _T_6144; // @[LoadQueue.scala 122:67:@11157.4]
  assign validEntriesInStoreQ_1 = _T_6113 ? _T_6135 : _T_6145; // @[LoadQueue.scala 121:91:@11158.4]
  assign _T_6149 = io_storeHead <= 4'h2; // @[LoadQueue.scala 122:18:@11160.4]
  assign _T_6151 = 4'h2 < io_storeTail; // @[LoadQueue.scala 122:36:@11161.4]
  assign _T_6152 = _T_6149 & _T_6151; // @[LoadQueue.scala 122:27:@11162.4]
  assign _T_6156 = io_storeTail <= 4'h2; // @[LoadQueue.scala 122:85:@11164.4]
  assign _T_6158 = 4'h2 < io_storeHead; // @[LoadQueue.scala 122:103:@11165.4]
  assign _T_6159 = _T_6156 & _T_6158; // @[LoadQueue.scala 122:94:@11166.4]
  assign _T_6161 = _T_6159 == 1'h0; // @[LoadQueue.scala 122:70:@11167.4]
  assign _T_6162 = _T_6120 & _T_6161; // @[LoadQueue.scala 122:67:@11168.4]
  assign validEntriesInStoreQ_2 = _T_6113 ? _T_6152 : _T_6162; // @[LoadQueue.scala 121:91:@11169.4]
  assign _T_6166 = io_storeHead <= 4'h3; // @[LoadQueue.scala 122:18:@11171.4]
  assign _T_6168 = 4'h3 < io_storeTail; // @[LoadQueue.scala 122:36:@11172.4]
  assign _T_6169 = _T_6166 & _T_6168; // @[LoadQueue.scala 122:27:@11173.4]
  assign _T_6173 = io_storeTail <= 4'h3; // @[LoadQueue.scala 122:85:@11175.4]
  assign _T_6175 = 4'h3 < io_storeHead; // @[LoadQueue.scala 122:103:@11176.4]
  assign _T_6176 = _T_6173 & _T_6175; // @[LoadQueue.scala 122:94:@11177.4]
  assign _T_6178 = _T_6176 == 1'h0; // @[LoadQueue.scala 122:70:@11178.4]
  assign _T_6179 = _T_6120 & _T_6178; // @[LoadQueue.scala 122:67:@11179.4]
  assign validEntriesInStoreQ_3 = _T_6113 ? _T_6169 : _T_6179; // @[LoadQueue.scala 121:91:@11180.4]
  assign _T_6183 = io_storeHead <= 4'h4; // @[LoadQueue.scala 122:18:@11182.4]
  assign _T_6185 = 4'h4 < io_storeTail; // @[LoadQueue.scala 122:36:@11183.4]
  assign _T_6186 = _T_6183 & _T_6185; // @[LoadQueue.scala 122:27:@11184.4]
  assign _T_6190 = io_storeTail <= 4'h4; // @[LoadQueue.scala 122:85:@11186.4]
  assign _T_6192 = 4'h4 < io_storeHead; // @[LoadQueue.scala 122:103:@11187.4]
  assign _T_6193 = _T_6190 & _T_6192; // @[LoadQueue.scala 122:94:@11188.4]
  assign _T_6195 = _T_6193 == 1'h0; // @[LoadQueue.scala 122:70:@11189.4]
  assign _T_6196 = _T_6120 & _T_6195; // @[LoadQueue.scala 122:67:@11190.4]
  assign validEntriesInStoreQ_4 = _T_6113 ? _T_6186 : _T_6196; // @[LoadQueue.scala 121:91:@11191.4]
  assign _T_6200 = io_storeHead <= 4'h5; // @[LoadQueue.scala 122:18:@11193.4]
  assign _T_6202 = 4'h5 < io_storeTail; // @[LoadQueue.scala 122:36:@11194.4]
  assign _T_6203 = _T_6200 & _T_6202; // @[LoadQueue.scala 122:27:@11195.4]
  assign _T_6207 = io_storeTail <= 4'h5; // @[LoadQueue.scala 122:85:@11197.4]
  assign _T_6209 = 4'h5 < io_storeHead; // @[LoadQueue.scala 122:103:@11198.4]
  assign _T_6210 = _T_6207 & _T_6209; // @[LoadQueue.scala 122:94:@11199.4]
  assign _T_6212 = _T_6210 == 1'h0; // @[LoadQueue.scala 122:70:@11200.4]
  assign _T_6213 = _T_6120 & _T_6212; // @[LoadQueue.scala 122:67:@11201.4]
  assign validEntriesInStoreQ_5 = _T_6113 ? _T_6203 : _T_6213; // @[LoadQueue.scala 121:91:@11202.4]
  assign _T_6217 = io_storeHead <= 4'h6; // @[LoadQueue.scala 122:18:@11204.4]
  assign _T_6219 = 4'h6 < io_storeTail; // @[LoadQueue.scala 122:36:@11205.4]
  assign _T_6220 = _T_6217 & _T_6219; // @[LoadQueue.scala 122:27:@11206.4]
  assign _T_6224 = io_storeTail <= 4'h6; // @[LoadQueue.scala 122:85:@11208.4]
  assign _T_6226 = 4'h6 < io_storeHead; // @[LoadQueue.scala 122:103:@11209.4]
  assign _T_6227 = _T_6224 & _T_6226; // @[LoadQueue.scala 122:94:@11210.4]
  assign _T_6229 = _T_6227 == 1'h0; // @[LoadQueue.scala 122:70:@11211.4]
  assign _T_6230 = _T_6120 & _T_6229; // @[LoadQueue.scala 122:67:@11212.4]
  assign validEntriesInStoreQ_6 = _T_6113 ? _T_6220 : _T_6230; // @[LoadQueue.scala 121:91:@11213.4]
  assign _T_6234 = io_storeHead <= 4'h7; // @[LoadQueue.scala 122:18:@11215.4]
  assign _T_6236 = 4'h7 < io_storeTail; // @[LoadQueue.scala 122:36:@11216.4]
  assign _T_6237 = _T_6234 & _T_6236; // @[LoadQueue.scala 122:27:@11217.4]
  assign _T_6241 = io_storeTail <= 4'h7; // @[LoadQueue.scala 122:85:@11219.4]
  assign _T_6243 = 4'h7 < io_storeHead; // @[LoadQueue.scala 122:103:@11220.4]
  assign _T_6244 = _T_6241 & _T_6243; // @[LoadQueue.scala 122:94:@11221.4]
  assign _T_6246 = _T_6244 == 1'h0; // @[LoadQueue.scala 122:70:@11222.4]
  assign _T_6247 = _T_6120 & _T_6246; // @[LoadQueue.scala 122:67:@11223.4]
  assign validEntriesInStoreQ_7 = _T_6113 ? _T_6237 : _T_6247; // @[LoadQueue.scala 121:91:@11224.4]
  assign _T_6251 = io_storeHead <= 4'h8; // @[LoadQueue.scala 122:18:@11226.4]
  assign _T_6253 = 4'h8 < io_storeTail; // @[LoadQueue.scala 122:36:@11227.4]
  assign _T_6254 = _T_6251 & _T_6253; // @[LoadQueue.scala 122:27:@11228.4]
  assign _T_6258 = io_storeTail <= 4'h8; // @[LoadQueue.scala 122:85:@11230.4]
  assign _T_6260 = 4'h8 < io_storeHead; // @[LoadQueue.scala 122:103:@11231.4]
  assign _T_6261 = _T_6258 & _T_6260; // @[LoadQueue.scala 122:94:@11232.4]
  assign _T_6263 = _T_6261 == 1'h0; // @[LoadQueue.scala 122:70:@11233.4]
  assign _T_6264 = _T_6120 & _T_6263; // @[LoadQueue.scala 122:67:@11234.4]
  assign validEntriesInStoreQ_8 = _T_6113 ? _T_6254 : _T_6264; // @[LoadQueue.scala 121:91:@11235.4]
  assign _T_6268 = io_storeHead <= 4'h9; // @[LoadQueue.scala 122:18:@11237.4]
  assign _T_6270 = 4'h9 < io_storeTail; // @[LoadQueue.scala 122:36:@11238.4]
  assign _T_6271 = _T_6268 & _T_6270; // @[LoadQueue.scala 122:27:@11239.4]
  assign _T_6275 = io_storeTail <= 4'h9; // @[LoadQueue.scala 122:85:@11241.4]
  assign _T_6277 = 4'h9 < io_storeHead; // @[LoadQueue.scala 122:103:@11242.4]
  assign _T_6278 = _T_6275 & _T_6277; // @[LoadQueue.scala 122:94:@11243.4]
  assign _T_6280 = _T_6278 == 1'h0; // @[LoadQueue.scala 122:70:@11244.4]
  assign _T_6281 = _T_6120 & _T_6280; // @[LoadQueue.scala 122:67:@11245.4]
  assign validEntriesInStoreQ_9 = _T_6113 ? _T_6271 : _T_6281; // @[LoadQueue.scala 121:91:@11246.4]
  assign _T_6285 = io_storeHead <= 4'ha; // @[LoadQueue.scala 122:18:@11248.4]
  assign _T_6287 = 4'ha < io_storeTail; // @[LoadQueue.scala 122:36:@11249.4]
  assign _T_6288 = _T_6285 & _T_6287; // @[LoadQueue.scala 122:27:@11250.4]
  assign _T_6292 = io_storeTail <= 4'ha; // @[LoadQueue.scala 122:85:@11252.4]
  assign _T_6294 = 4'ha < io_storeHead; // @[LoadQueue.scala 122:103:@11253.4]
  assign _T_6295 = _T_6292 & _T_6294; // @[LoadQueue.scala 122:94:@11254.4]
  assign _T_6297 = _T_6295 == 1'h0; // @[LoadQueue.scala 122:70:@11255.4]
  assign _T_6298 = _T_6120 & _T_6297; // @[LoadQueue.scala 122:67:@11256.4]
  assign validEntriesInStoreQ_10 = _T_6113 ? _T_6288 : _T_6298; // @[LoadQueue.scala 121:91:@11257.4]
  assign _T_6302 = io_storeHead <= 4'hb; // @[LoadQueue.scala 122:18:@11259.4]
  assign _T_6304 = 4'hb < io_storeTail; // @[LoadQueue.scala 122:36:@11260.4]
  assign _T_6305 = _T_6302 & _T_6304; // @[LoadQueue.scala 122:27:@11261.4]
  assign _T_6309 = io_storeTail <= 4'hb; // @[LoadQueue.scala 122:85:@11263.4]
  assign _T_6311 = 4'hb < io_storeHead; // @[LoadQueue.scala 122:103:@11264.4]
  assign _T_6312 = _T_6309 & _T_6311; // @[LoadQueue.scala 122:94:@11265.4]
  assign _T_6314 = _T_6312 == 1'h0; // @[LoadQueue.scala 122:70:@11266.4]
  assign _T_6315 = _T_6120 & _T_6314; // @[LoadQueue.scala 122:67:@11267.4]
  assign validEntriesInStoreQ_11 = _T_6113 ? _T_6305 : _T_6315; // @[LoadQueue.scala 121:91:@11268.4]
  assign _T_6319 = io_storeHead <= 4'hc; // @[LoadQueue.scala 122:18:@11270.4]
  assign _T_6321 = 4'hc < io_storeTail; // @[LoadQueue.scala 122:36:@11271.4]
  assign _T_6322 = _T_6319 & _T_6321; // @[LoadQueue.scala 122:27:@11272.4]
  assign _T_6326 = io_storeTail <= 4'hc; // @[LoadQueue.scala 122:85:@11274.4]
  assign _T_6328 = 4'hc < io_storeHead; // @[LoadQueue.scala 122:103:@11275.4]
  assign _T_6329 = _T_6326 & _T_6328; // @[LoadQueue.scala 122:94:@11276.4]
  assign _T_6331 = _T_6329 == 1'h0; // @[LoadQueue.scala 122:70:@11277.4]
  assign _T_6332 = _T_6120 & _T_6331; // @[LoadQueue.scala 122:67:@11278.4]
  assign validEntriesInStoreQ_12 = _T_6113 ? _T_6322 : _T_6332; // @[LoadQueue.scala 121:91:@11279.4]
  assign _T_6336 = io_storeHead <= 4'hd; // @[LoadQueue.scala 122:18:@11281.4]
  assign _T_6338 = 4'hd < io_storeTail; // @[LoadQueue.scala 122:36:@11282.4]
  assign _T_6339 = _T_6336 & _T_6338; // @[LoadQueue.scala 122:27:@11283.4]
  assign _T_6343 = io_storeTail <= 4'hd; // @[LoadQueue.scala 122:85:@11285.4]
  assign _T_6345 = 4'hd < io_storeHead; // @[LoadQueue.scala 122:103:@11286.4]
  assign _T_6346 = _T_6343 & _T_6345; // @[LoadQueue.scala 122:94:@11287.4]
  assign _T_6348 = _T_6346 == 1'h0; // @[LoadQueue.scala 122:70:@11288.4]
  assign _T_6349 = _T_6120 & _T_6348; // @[LoadQueue.scala 122:67:@11289.4]
  assign validEntriesInStoreQ_13 = _T_6113 ? _T_6339 : _T_6349; // @[LoadQueue.scala 121:91:@11290.4]
  assign _T_6353 = io_storeHead <= 4'he; // @[LoadQueue.scala 122:18:@11292.4]
  assign _T_6355 = 4'he < io_storeTail; // @[LoadQueue.scala 122:36:@11293.4]
  assign _T_6356 = _T_6353 & _T_6355; // @[LoadQueue.scala 122:27:@11294.4]
  assign _T_6360 = io_storeTail <= 4'he; // @[LoadQueue.scala 122:85:@11296.4]
  assign _T_6362 = 4'he < io_storeHead; // @[LoadQueue.scala 122:103:@11297.4]
  assign _T_6363 = _T_6360 & _T_6362; // @[LoadQueue.scala 122:94:@11298.4]
  assign _T_6365 = _T_6363 == 1'h0; // @[LoadQueue.scala 122:70:@11299.4]
  assign _T_6366 = _T_6120 & _T_6365; // @[LoadQueue.scala 122:67:@11300.4]
  assign validEntriesInStoreQ_14 = _T_6113 ? _T_6356 : _T_6366; // @[LoadQueue.scala 121:91:@11301.4]
  assign validEntriesInStoreQ_15 = _T_6113 ? 1'h0 : _T_6120; // @[LoadQueue.scala 121:91:@11312.4]
  assign storesToCheck_0_0 = _T_2228 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11339.4]
  assign _T_7654 = 4'h1 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11342.4]
  assign _T_7655 = _T_6132 & _T_7654; // @[LoadQueue.scala 131:72:@11343.4]
  assign _T_7657 = offsetQ_0 < 4'h1; // @[LoadQueue.scala 132:33:@11344.4]
  assign _T_7660 = _T_7657 & _T_6141; // @[LoadQueue.scala 132:41:@11346.4]
  assign _T_7662 = _T_7660 == 1'h0; // @[LoadQueue.scala 132:9:@11347.4]
  assign storesToCheck_0_1 = _T_2228 ? _T_7655 : _T_7662; // @[LoadQueue.scala 131:10:@11348.4]
  assign _T_7668 = 4'h2 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11351.4]
  assign _T_7669 = _T_6149 & _T_7668; // @[LoadQueue.scala 131:72:@11352.4]
  assign _T_7671 = offsetQ_0 < 4'h2; // @[LoadQueue.scala 132:33:@11353.4]
  assign _T_7674 = _T_7671 & _T_6158; // @[LoadQueue.scala 132:41:@11355.4]
  assign _T_7676 = _T_7674 == 1'h0; // @[LoadQueue.scala 132:9:@11356.4]
  assign storesToCheck_0_2 = _T_2228 ? _T_7669 : _T_7676; // @[LoadQueue.scala 131:10:@11357.4]
  assign _T_7682 = 4'h3 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11360.4]
  assign _T_7683 = _T_6166 & _T_7682; // @[LoadQueue.scala 131:72:@11361.4]
  assign _T_7685 = offsetQ_0 < 4'h3; // @[LoadQueue.scala 132:33:@11362.4]
  assign _T_7688 = _T_7685 & _T_6175; // @[LoadQueue.scala 132:41:@11364.4]
  assign _T_7690 = _T_7688 == 1'h0; // @[LoadQueue.scala 132:9:@11365.4]
  assign storesToCheck_0_3 = _T_2228 ? _T_7683 : _T_7690; // @[LoadQueue.scala 131:10:@11366.4]
  assign _T_7696 = 4'h4 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11369.4]
  assign _T_7697 = _T_6183 & _T_7696; // @[LoadQueue.scala 131:72:@11370.4]
  assign _T_7699 = offsetQ_0 < 4'h4; // @[LoadQueue.scala 132:33:@11371.4]
  assign _T_7702 = _T_7699 & _T_6192; // @[LoadQueue.scala 132:41:@11373.4]
  assign _T_7704 = _T_7702 == 1'h0; // @[LoadQueue.scala 132:9:@11374.4]
  assign storesToCheck_0_4 = _T_2228 ? _T_7697 : _T_7704; // @[LoadQueue.scala 131:10:@11375.4]
  assign _T_7710 = 4'h5 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11378.4]
  assign _T_7711 = _T_6200 & _T_7710; // @[LoadQueue.scala 131:72:@11379.4]
  assign _T_7713 = offsetQ_0 < 4'h5; // @[LoadQueue.scala 132:33:@11380.4]
  assign _T_7716 = _T_7713 & _T_6209; // @[LoadQueue.scala 132:41:@11382.4]
  assign _T_7718 = _T_7716 == 1'h0; // @[LoadQueue.scala 132:9:@11383.4]
  assign storesToCheck_0_5 = _T_2228 ? _T_7711 : _T_7718; // @[LoadQueue.scala 131:10:@11384.4]
  assign _T_7724 = 4'h6 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11387.4]
  assign _T_7725 = _T_6217 & _T_7724; // @[LoadQueue.scala 131:72:@11388.4]
  assign _T_7727 = offsetQ_0 < 4'h6; // @[LoadQueue.scala 132:33:@11389.4]
  assign _T_7730 = _T_7727 & _T_6226; // @[LoadQueue.scala 132:41:@11391.4]
  assign _T_7732 = _T_7730 == 1'h0; // @[LoadQueue.scala 132:9:@11392.4]
  assign storesToCheck_0_6 = _T_2228 ? _T_7725 : _T_7732; // @[LoadQueue.scala 131:10:@11393.4]
  assign _T_7738 = 4'h7 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11396.4]
  assign _T_7739 = _T_6234 & _T_7738; // @[LoadQueue.scala 131:72:@11397.4]
  assign _T_7741 = offsetQ_0 < 4'h7; // @[LoadQueue.scala 132:33:@11398.4]
  assign _T_7744 = _T_7741 & _T_6243; // @[LoadQueue.scala 132:41:@11400.4]
  assign _T_7746 = _T_7744 == 1'h0; // @[LoadQueue.scala 132:9:@11401.4]
  assign storesToCheck_0_7 = _T_2228 ? _T_7739 : _T_7746; // @[LoadQueue.scala 131:10:@11402.4]
  assign _T_7752 = 4'h8 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11405.4]
  assign _T_7753 = _T_6251 & _T_7752; // @[LoadQueue.scala 131:72:@11406.4]
  assign _T_7755 = offsetQ_0 < 4'h8; // @[LoadQueue.scala 132:33:@11407.4]
  assign _T_7758 = _T_7755 & _T_6260; // @[LoadQueue.scala 132:41:@11409.4]
  assign _T_7760 = _T_7758 == 1'h0; // @[LoadQueue.scala 132:9:@11410.4]
  assign storesToCheck_0_8 = _T_2228 ? _T_7753 : _T_7760; // @[LoadQueue.scala 131:10:@11411.4]
  assign _T_7766 = 4'h9 <= offsetQ_0; // @[LoadQueue.scala 131:81:@11414.4]
  assign _T_7767 = _T_6268 & _T_7766; // @[LoadQueue.scala 131:72:@11415.4]
  assign _T_7769 = offsetQ_0 < 4'h9; // @[LoadQueue.scala 132:33:@11416.4]
  assign _T_7772 = _T_7769 & _T_6277; // @[LoadQueue.scala 132:41:@11418.4]
  assign _T_7774 = _T_7772 == 1'h0; // @[LoadQueue.scala 132:9:@11419.4]
  assign storesToCheck_0_9 = _T_2228 ? _T_7767 : _T_7774; // @[LoadQueue.scala 131:10:@11420.4]
  assign _T_7780 = 4'ha <= offsetQ_0; // @[LoadQueue.scala 131:81:@11423.4]
  assign _T_7781 = _T_6285 & _T_7780; // @[LoadQueue.scala 131:72:@11424.4]
  assign _T_7783 = offsetQ_0 < 4'ha; // @[LoadQueue.scala 132:33:@11425.4]
  assign _T_7786 = _T_7783 & _T_6294; // @[LoadQueue.scala 132:41:@11427.4]
  assign _T_7788 = _T_7786 == 1'h0; // @[LoadQueue.scala 132:9:@11428.4]
  assign storesToCheck_0_10 = _T_2228 ? _T_7781 : _T_7788; // @[LoadQueue.scala 131:10:@11429.4]
  assign _T_7794 = 4'hb <= offsetQ_0; // @[LoadQueue.scala 131:81:@11432.4]
  assign _T_7795 = _T_6302 & _T_7794; // @[LoadQueue.scala 131:72:@11433.4]
  assign _T_7797 = offsetQ_0 < 4'hb; // @[LoadQueue.scala 132:33:@11434.4]
  assign _T_7800 = _T_7797 & _T_6311; // @[LoadQueue.scala 132:41:@11436.4]
  assign _T_7802 = _T_7800 == 1'h0; // @[LoadQueue.scala 132:9:@11437.4]
  assign storesToCheck_0_11 = _T_2228 ? _T_7795 : _T_7802; // @[LoadQueue.scala 131:10:@11438.4]
  assign _T_7808 = 4'hc <= offsetQ_0; // @[LoadQueue.scala 131:81:@11441.4]
  assign _T_7809 = _T_6319 & _T_7808; // @[LoadQueue.scala 131:72:@11442.4]
  assign _T_7811 = offsetQ_0 < 4'hc; // @[LoadQueue.scala 132:33:@11443.4]
  assign _T_7814 = _T_7811 & _T_6328; // @[LoadQueue.scala 132:41:@11445.4]
  assign _T_7816 = _T_7814 == 1'h0; // @[LoadQueue.scala 132:9:@11446.4]
  assign storesToCheck_0_12 = _T_2228 ? _T_7809 : _T_7816; // @[LoadQueue.scala 131:10:@11447.4]
  assign _T_7822 = 4'hd <= offsetQ_0; // @[LoadQueue.scala 131:81:@11450.4]
  assign _T_7823 = _T_6336 & _T_7822; // @[LoadQueue.scala 131:72:@11451.4]
  assign _T_7825 = offsetQ_0 < 4'hd; // @[LoadQueue.scala 132:33:@11452.4]
  assign _T_7828 = _T_7825 & _T_6345; // @[LoadQueue.scala 132:41:@11454.4]
  assign _T_7830 = _T_7828 == 1'h0; // @[LoadQueue.scala 132:9:@11455.4]
  assign storesToCheck_0_13 = _T_2228 ? _T_7823 : _T_7830; // @[LoadQueue.scala 131:10:@11456.4]
  assign _T_7836 = 4'he <= offsetQ_0; // @[LoadQueue.scala 131:81:@11459.4]
  assign _T_7837 = _T_6353 & _T_7836; // @[LoadQueue.scala 131:72:@11460.4]
  assign _T_7839 = offsetQ_0 < 4'he; // @[LoadQueue.scala 132:33:@11461.4]
  assign _T_7842 = _T_7839 & _T_6362; // @[LoadQueue.scala 132:41:@11463.4]
  assign _T_7844 = _T_7842 == 1'h0; // @[LoadQueue.scala 132:9:@11464.4]
  assign storesToCheck_0_14 = _T_2228 ? _T_7837 : _T_7844; // @[LoadQueue.scala 131:10:@11465.4]
  assign _T_7850 = 4'hf <= offsetQ_0; // @[LoadQueue.scala 131:81:@11468.4]
  assign storesToCheck_0_15 = _T_2228 ? _T_7850 : 1'h1; // @[LoadQueue.scala 131:10:@11474.4]
  assign storesToCheck_1_0 = _T_2258 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11516.4]
  assign _T_7900 = 4'h1 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11519.4]
  assign _T_7901 = _T_6132 & _T_7900; // @[LoadQueue.scala 131:72:@11520.4]
  assign _T_7903 = offsetQ_1 < 4'h1; // @[LoadQueue.scala 132:33:@11521.4]
  assign _T_7906 = _T_7903 & _T_6141; // @[LoadQueue.scala 132:41:@11523.4]
  assign _T_7908 = _T_7906 == 1'h0; // @[LoadQueue.scala 132:9:@11524.4]
  assign storesToCheck_1_1 = _T_2258 ? _T_7901 : _T_7908; // @[LoadQueue.scala 131:10:@11525.4]
  assign _T_7914 = 4'h2 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11528.4]
  assign _T_7915 = _T_6149 & _T_7914; // @[LoadQueue.scala 131:72:@11529.4]
  assign _T_7917 = offsetQ_1 < 4'h2; // @[LoadQueue.scala 132:33:@11530.4]
  assign _T_7920 = _T_7917 & _T_6158; // @[LoadQueue.scala 132:41:@11532.4]
  assign _T_7922 = _T_7920 == 1'h0; // @[LoadQueue.scala 132:9:@11533.4]
  assign storesToCheck_1_2 = _T_2258 ? _T_7915 : _T_7922; // @[LoadQueue.scala 131:10:@11534.4]
  assign _T_7928 = 4'h3 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11537.4]
  assign _T_7929 = _T_6166 & _T_7928; // @[LoadQueue.scala 131:72:@11538.4]
  assign _T_7931 = offsetQ_1 < 4'h3; // @[LoadQueue.scala 132:33:@11539.4]
  assign _T_7934 = _T_7931 & _T_6175; // @[LoadQueue.scala 132:41:@11541.4]
  assign _T_7936 = _T_7934 == 1'h0; // @[LoadQueue.scala 132:9:@11542.4]
  assign storesToCheck_1_3 = _T_2258 ? _T_7929 : _T_7936; // @[LoadQueue.scala 131:10:@11543.4]
  assign _T_7942 = 4'h4 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11546.4]
  assign _T_7943 = _T_6183 & _T_7942; // @[LoadQueue.scala 131:72:@11547.4]
  assign _T_7945 = offsetQ_1 < 4'h4; // @[LoadQueue.scala 132:33:@11548.4]
  assign _T_7948 = _T_7945 & _T_6192; // @[LoadQueue.scala 132:41:@11550.4]
  assign _T_7950 = _T_7948 == 1'h0; // @[LoadQueue.scala 132:9:@11551.4]
  assign storesToCheck_1_4 = _T_2258 ? _T_7943 : _T_7950; // @[LoadQueue.scala 131:10:@11552.4]
  assign _T_7956 = 4'h5 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11555.4]
  assign _T_7957 = _T_6200 & _T_7956; // @[LoadQueue.scala 131:72:@11556.4]
  assign _T_7959 = offsetQ_1 < 4'h5; // @[LoadQueue.scala 132:33:@11557.4]
  assign _T_7962 = _T_7959 & _T_6209; // @[LoadQueue.scala 132:41:@11559.4]
  assign _T_7964 = _T_7962 == 1'h0; // @[LoadQueue.scala 132:9:@11560.4]
  assign storesToCheck_1_5 = _T_2258 ? _T_7957 : _T_7964; // @[LoadQueue.scala 131:10:@11561.4]
  assign _T_7970 = 4'h6 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11564.4]
  assign _T_7971 = _T_6217 & _T_7970; // @[LoadQueue.scala 131:72:@11565.4]
  assign _T_7973 = offsetQ_1 < 4'h6; // @[LoadQueue.scala 132:33:@11566.4]
  assign _T_7976 = _T_7973 & _T_6226; // @[LoadQueue.scala 132:41:@11568.4]
  assign _T_7978 = _T_7976 == 1'h0; // @[LoadQueue.scala 132:9:@11569.4]
  assign storesToCheck_1_6 = _T_2258 ? _T_7971 : _T_7978; // @[LoadQueue.scala 131:10:@11570.4]
  assign _T_7984 = 4'h7 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11573.4]
  assign _T_7985 = _T_6234 & _T_7984; // @[LoadQueue.scala 131:72:@11574.4]
  assign _T_7987 = offsetQ_1 < 4'h7; // @[LoadQueue.scala 132:33:@11575.4]
  assign _T_7990 = _T_7987 & _T_6243; // @[LoadQueue.scala 132:41:@11577.4]
  assign _T_7992 = _T_7990 == 1'h0; // @[LoadQueue.scala 132:9:@11578.4]
  assign storesToCheck_1_7 = _T_2258 ? _T_7985 : _T_7992; // @[LoadQueue.scala 131:10:@11579.4]
  assign _T_7998 = 4'h8 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11582.4]
  assign _T_7999 = _T_6251 & _T_7998; // @[LoadQueue.scala 131:72:@11583.4]
  assign _T_8001 = offsetQ_1 < 4'h8; // @[LoadQueue.scala 132:33:@11584.4]
  assign _T_8004 = _T_8001 & _T_6260; // @[LoadQueue.scala 132:41:@11586.4]
  assign _T_8006 = _T_8004 == 1'h0; // @[LoadQueue.scala 132:9:@11587.4]
  assign storesToCheck_1_8 = _T_2258 ? _T_7999 : _T_8006; // @[LoadQueue.scala 131:10:@11588.4]
  assign _T_8012 = 4'h9 <= offsetQ_1; // @[LoadQueue.scala 131:81:@11591.4]
  assign _T_8013 = _T_6268 & _T_8012; // @[LoadQueue.scala 131:72:@11592.4]
  assign _T_8015 = offsetQ_1 < 4'h9; // @[LoadQueue.scala 132:33:@11593.4]
  assign _T_8018 = _T_8015 & _T_6277; // @[LoadQueue.scala 132:41:@11595.4]
  assign _T_8020 = _T_8018 == 1'h0; // @[LoadQueue.scala 132:9:@11596.4]
  assign storesToCheck_1_9 = _T_2258 ? _T_8013 : _T_8020; // @[LoadQueue.scala 131:10:@11597.4]
  assign _T_8026 = 4'ha <= offsetQ_1; // @[LoadQueue.scala 131:81:@11600.4]
  assign _T_8027 = _T_6285 & _T_8026; // @[LoadQueue.scala 131:72:@11601.4]
  assign _T_8029 = offsetQ_1 < 4'ha; // @[LoadQueue.scala 132:33:@11602.4]
  assign _T_8032 = _T_8029 & _T_6294; // @[LoadQueue.scala 132:41:@11604.4]
  assign _T_8034 = _T_8032 == 1'h0; // @[LoadQueue.scala 132:9:@11605.4]
  assign storesToCheck_1_10 = _T_2258 ? _T_8027 : _T_8034; // @[LoadQueue.scala 131:10:@11606.4]
  assign _T_8040 = 4'hb <= offsetQ_1; // @[LoadQueue.scala 131:81:@11609.4]
  assign _T_8041 = _T_6302 & _T_8040; // @[LoadQueue.scala 131:72:@11610.4]
  assign _T_8043 = offsetQ_1 < 4'hb; // @[LoadQueue.scala 132:33:@11611.4]
  assign _T_8046 = _T_8043 & _T_6311; // @[LoadQueue.scala 132:41:@11613.4]
  assign _T_8048 = _T_8046 == 1'h0; // @[LoadQueue.scala 132:9:@11614.4]
  assign storesToCheck_1_11 = _T_2258 ? _T_8041 : _T_8048; // @[LoadQueue.scala 131:10:@11615.4]
  assign _T_8054 = 4'hc <= offsetQ_1; // @[LoadQueue.scala 131:81:@11618.4]
  assign _T_8055 = _T_6319 & _T_8054; // @[LoadQueue.scala 131:72:@11619.4]
  assign _T_8057 = offsetQ_1 < 4'hc; // @[LoadQueue.scala 132:33:@11620.4]
  assign _T_8060 = _T_8057 & _T_6328; // @[LoadQueue.scala 132:41:@11622.4]
  assign _T_8062 = _T_8060 == 1'h0; // @[LoadQueue.scala 132:9:@11623.4]
  assign storesToCheck_1_12 = _T_2258 ? _T_8055 : _T_8062; // @[LoadQueue.scala 131:10:@11624.4]
  assign _T_8068 = 4'hd <= offsetQ_1; // @[LoadQueue.scala 131:81:@11627.4]
  assign _T_8069 = _T_6336 & _T_8068; // @[LoadQueue.scala 131:72:@11628.4]
  assign _T_8071 = offsetQ_1 < 4'hd; // @[LoadQueue.scala 132:33:@11629.4]
  assign _T_8074 = _T_8071 & _T_6345; // @[LoadQueue.scala 132:41:@11631.4]
  assign _T_8076 = _T_8074 == 1'h0; // @[LoadQueue.scala 132:9:@11632.4]
  assign storesToCheck_1_13 = _T_2258 ? _T_8069 : _T_8076; // @[LoadQueue.scala 131:10:@11633.4]
  assign _T_8082 = 4'he <= offsetQ_1; // @[LoadQueue.scala 131:81:@11636.4]
  assign _T_8083 = _T_6353 & _T_8082; // @[LoadQueue.scala 131:72:@11637.4]
  assign _T_8085 = offsetQ_1 < 4'he; // @[LoadQueue.scala 132:33:@11638.4]
  assign _T_8088 = _T_8085 & _T_6362; // @[LoadQueue.scala 132:41:@11640.4]
  assign _T_8090 = _T_8088 == 1'h0; // @[LoadQueue.scala 132:9:@11641.4]
  assign storesToCheck_1_14 = _T_2258 ? _T_8083 : _T_8090; // @[LoadQueue.scala 131:10:@11642.4]
  assign _T_8096 = 4'hf <= offsetQ_1; // @[LoadQueue.scala 131:81:@11645.4]
  assign storesToCheck_1_15 = _T_2258 ? _T_8096 : 1'h1; // @[LoadQueue.scala 131:10:@11651.4]
  assign storesToCheck_2_0 = _T_2288 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11693.4]
  assign _T_8146 = 4'h1 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11696.4]
  assign _T_8147 = _T_6132 & _T_8146; // @[LoadQueue.scala 131:72:@11697.4]
  assign _T_8149 = offsetQ_2 < 4'h1; // @[LoadQueue.scala 132:33:@11698.4]
  assign _T_8152 = _T_8149 & _T_6141; // @[LoadQueue.scala 132:41:@11700.4]
  assign _T_8154 = _T_8152 == 1'h0; // @[LoadQueue.scala 132:9:@11701.4]
  assign storesToCheck_2_1 = _T_2288 ? _T_8147 : _T_8154; // @[LoadQueue.scala 131:10:@11702.4]
  assign _T_8160 = 4'h2 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11705.4]
  assign _T_8161 = _T_6149 & _T_8160; // @[LoadQueue.scala 131:72:@11706.4]
  assign _T_8163 = offsetQ_2 < 4'h2; // @[LoadQueue.scala 132:33:@11707.4]
  assign _T_8166 = _T_8163 & _T_6158; // @[LoadQueue.scala 132:41:@11709.4]
  assign _T_8168 = _T_8166 == 1'h0; // @[LoadQueue.scala 132:9:@11710.4]
  assign storesToCheck_2_2 = _T_2288 ? _T_8161 : _T_8168; // @[LoadQueue.scala 131:10:@11711.4]
  assign _T_8174 = 4'h3 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11714.4]
  assign _T_8175 = _T_6166 & _T_8174; // @[LoadQueue.scala 131:72:@11715.4]
  assign _T_8177 = offsetQ_2 < 4'h3; // @[LoadQueue.scala 132:33:@11716.4]
  assign _T_8180 = _T_8177 & _T_6175; // @[LoadQueue.scala 132:41:@11718.4]
  assign _T_8182 = _T_8180 == 1'h0; // @[LoadQueue.scala 132:9:@11719.4]
  assign storesToCheck_2_3 = _T_2288 ? _T_8175 : _T_8182; // @[LoadQueue.scala 131:10:@11720.4]
  assign _T_8188 = 4'h4 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11723.4]
  assign _T_8189 = _T_6183 & _T_8188; // @[LoadQueue.scala 131:72:@11724.4]
  assign _T_8191 = offsetQ_2 < 4'h4; // @[LoadQueue.scala 132:33:@11725.4]
  assign _T_8194 = _T_8191 & _T_6192; // @[LoadQueue.scala 132:41:@11727.4]
  assign _T_8196 = _T_8194 == 1'h0; // @[LoadQueue.scala 132:9:@11728.4]
  assign storesToCheck_2_4 = _T_2288 ? _T_8189 : _T_8196; // @[LoadQueue.scala 131:10:@11729.4]
  assign _T_8202 = 4'h5 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11732.4]
  assign _T_8203 = _T_6200 & _T_8202; // @[LoadQueue.scala 131:72:@11733.4]
  assign _T_8205 = offsetQ_2 < 4'h5; // @[LoadQueue.scala 132:33:@11734.4]
  assign _T_8208 = _T_8205 & _T_6209; // @[LoadQueue.scala 132:41:@11736.4]
  assign _T_8210 = _T_8208 == 1'h0; // @[LoadQueue.scala 132:9:@11737.4]
  assign storesToCheck_2_5 = _T_2288 ? _T_8203 : _T_8210; // @[LoadQueue.scala 131:10:@11738.4]
  assign _T_8216 = 4'h6 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11741.4]
  assign _T_8217 = _T_6217 & _T_8216; // @[LoadQueue.scala 131:72:@11742.4]
  assign _T_8219 = offsetQ_2 < 4'h6; // @[LoadQueue.scala 132:33:@11743.4]
  assign _T_8222 = _T_8219 & _T_6226; // @[LoadQueue.scala 132:41:@11745.4]
  assign _T_8224 = _T_8222 == 1'h0; // @[LoadQueue.scala 132:9:@11746.4]
  assign storesToCheck_2_6 = _T_2288 ? _T_8217 : _T_8224; // @[LoadQueue.scala 131:10:@11747.4]
  assign _T_8230 = 4'h7 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11750.4]
  assign _T_8231 = _T_6234 & _T_8230; // @[LoadQueue.scala 131:72:@11751.4]
  assign _T_8233 = offsetQ_2 < 4'h7; // @[LoadQueue.scala 132:33:@11752.4]
  assign _T_8236 = _T_8233 & _T_6243; // @[LoadQueue.scala 132:41:@11754.4]
  assign _T_8238 = _T_8236 == 1'h0; // @[LoadQueue.scala 132:9:@11755.4]
  assign storesToCheck_2_7 = _T_2288 ? _T_8231 : _T_8238; // @[LoadQueue.scala 131:10:@11756.4]
  assign _T_8244 = 4'h8 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11759.4]
  assign _T_8245 = _T_6251 & _T_8244; // @[LoadQueue.scala 131:72:@11760.4]
  assign _T_8247 = offsetQ_2 < 4'h8; // @[LoadQueue.scala 132:33:@11761.4]
  assign _T_8250 = _T_8247 & _T_6260; // @[LoadQueue.scala 132:41:@11763.4]
  assign _T_8252 = _T_8250 == 1'h0; // @[LoadQueue.scala 132:9:@11764.4]
  assign storesToCheck_2_8 = _T_2288 ? _T_8245 : _T_8252; // @[LoadQueue.scala 131:10:@11765.4]
  assign _T_8258 = 4'h9 <= offsetQ_2; // @[LoadQueue.scala 131:81:@11768.4]
  assign _T_8259 = _T_6268 & _T_8258; // @[LoadQueue.scala 131:72:@11769.4]
  assign _T_8261 = offsetQ_2 < 4'h9; // @[LoadQueue.scala 132:33:@11770.4]
  assign _T_8264 = _T_8261 & _T_6277; // @[LoadQueue.scala 132:41:@11772.4]
  assign _T_8266 = _T_8264 == 1'h0; // @[LoadQueue.scala 132:9:@11773.4]
  assign storesToCheck_2_9 = _T_2288 ? _T_8259 : _T_8266; // @[LoadQueue.scala 131:10:@11774.4]
  assign _T_8272 = 4'ha <= offsetQ_2; // @[LoadQueue.scala 131:81:@11777.4]
  assign _T_8273 = _T_6285 & _T_8272; // @[LoadQueue.scala 131:72:@11778.4]
  assign _T_8275 = offsetQ_2 < 4'ha; // @[LoadQueue.scala 132:33:@11779.4]
  assign _T_8278 = _T_8275 & _T_6294; // @[LoadQueue.scala 132:41:@11781.4]
  assign _T_8280 = _T_8278 == 1'h0; // @[LoadQueue.scala 132:9:@11782.4]
  assign storesToCheck_2_10 = _T_2288 ? _T_8273 : _T_8280; // @[LoadQueue.scala 131:10:@11783.4]
  assign _T_8286 = 4'hb <= offsetQ_2; // @[LoadQueue.scala 131:81:@11786.4]
  assign _T_8287 = _T_6302 & _T_8286; // @[LoadQueue.scala 131:72:@11787.4]
  assign _T_8289 = offsetQ_2 < 4'hb; // @[LoadQueue.scala 132:33:@11788.4]
  assign _T_8292 = _T_8289 & _T_6311; // @[LoadQueue.scala 132:41:@11790.4]
  assign _T_8294 = _T_8292 == 1'h0; // @[LoadQueue.scala 132:9:@11791.4]
  assign storesToCheck_2_11 = _T_2288 ? _T_8287 : _T_8294; // @[LoadQueue.scala 131:10:@11792.4]
  assign _T_8300 = 4'hc <= offsetQ_2; // @[LoadQueue.scala 131:81:@11795.4]
  assign _T_8301 = _T_6319 & _T_8300; // @[LoadQueue.scala 131:72:@11796.4]
  assign _T_8303 = offsetQ_2 < 4'hc; // @[LoadQueue.scala 132:33:@11797.4]
  assign _T_8306 = _T_8303 & _T_6328; // @[LoadQueue.scala 132:41:@11799.4]
  assign _T_8308 = _T_8306 == 1'h0; // @[LoadQueue.scala 132:9:@11800.4]
  assign storesToCheck_2_12 = _T_2288 ? _T_8301 : _T_8308; // @[LoadQueue.scala 131:10:@11801.4]
  assign _T_8314 = 4'hd <= offsetQ_2; // @[LoadQueue.scala 131:81:@11804.4]
  assign _T_8315 = _T_6336 & _T_8314; // @[LoadQueue.scala 131:72:@11805.4]
  assign _T_8317 = offsetQ_2 < 4'hd; // @[LoadQueue.scala 132:33:@11806.4]
  assign _T_8320 = _T_8317 & _T_6345; // @[LoadQueue.scala 132:41:@11808.4]
  assign _T_8322 = _T_8320 == 1'h0; // @[LoadQueue.scala 132:9:@11809.4]
  assign storesToCheck_2_13 = _T_2288 ? _T_8315 : _T_8322; // @[LoadQueue.scala 131:10:@11810.4]
  assign _T_8328 = 4'he <= offsetQ_2; // @[LoadQueue.scala 131:81:@11813.4]
  assign _T_8329 = _T_6353 & _T_8328; // @[LoadQueue.scala 131:72:@11814.4]
  assign _T_8331 = offsetQ_2 < 4'he; // @[LoadQueue.scala 132:33:@11815.4]
  assign _T_8334 = _T_8331 & _T_6362; // @[LoadQueue.scala 132:41:@11817.4]
  assign _T_8336 = _T_8334 == 1'h0; // @[LoadQueue.scala 132:9:@11818.4]
  assign storesToCheck_2_14 = _T_2288 ? _T_8329 : _T_8336; // @[LoadQueue.scala 131:10:@11819.4]
  assign _T_8342 = 4'hf <= offsetQ_2; // @[LoadQueue.scala 131:81:@11822.4]
  assign storesToCheck_2_15 = _T_2288 ? _T_8342 : 1'h1; // @[LoadQueue.scala 131:10:@11828.4]
  assign storesToCheck_3_0 = _T_2318 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11870.4]
  assign _T_8392 = 4'h1 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11873.4]
  assign _T_8393 = _T_6132 & _T_8392; // @[LoadQueue.scala 131:72:@11874.4]
  assign _T_8395 = offsetQ_3 < 4'h1; // @[LoadQueue.scala 132:33:@11875.4]
  assign _T_8398 = _T_8395 & _T_6141; // @[LoadQueue.scala 132:41:@11877.4]
  assign _T_8400 = _T_8398 == 1'h0; // @[LoadQueue.scala 132:9:@11878.4]
  assign storesToCheck_3_1 = _T_2318 ? _T_8393 : _T_8400; // @[LoadQueue.scala 131:10:@11879.4]
  assign _T_8406 = 4'h2 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11882.4]
  assign _T_8407 = _T_6149 & _T_8406; // @[LoadQueue.scala 131:72:@11883.4]
  assign _T_8409 = offsetQ_3 < 4'h2; // @[LoadQueue.scala 132:33:@11884.4]
  assign _T_8412 = _T_8409 & _T_6158; // @[LoadQueue.scala 132:41:@11886.4]
  assign _T_8414 = _T_8412 == 1'h0; // @[LoadQueue.scala 132:9:@11887.4]
  assign storesToCheck_3_2 = _T_2318 ? _T_8407 : _T_8414; // @[LoadQueue.scala 131:10:@11888.4]
  assign _T_8420 = 4'h3 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11891.4]
  assign _T_8421 = _T_6166 & _T_8420; // @[LoadQueue.scala 131:72:@11892.4]
  assign _T_8423 = offsetQ_3 < 4'h3; // @[LoadQueue.scala 132:33:@11893.4]
  assign _T_8426 = _T_8423 & _T_6175; // @[LoadQueue.scala 132:41:@11895.4]
  assign _T_8428 = _T_8426 == 1'h0; // @[LoadQueue.scala 132:9:@11896.4]
  assign storesToCheck_3_3 = _T_2318 ? _T_8421 : _T_8428; // @[LoadQueue.scala 131:10:@11897.4]
  assign _T_8434 = 4'h4 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11900.4]
  assign _T_8435 = _T_6183 & _T_8434; // @[LoadQueue.scala 131:72:@11901.4]
  assign _T_8437 = offsetQ_3 < 4'h4; // @[LoadQueue.scala 132:33:@11902.4]
  assign _T_8440 = _T_8437 & _T_6192; // @[LoadQueue.scala 132:41:@11904.4]
  assign _T_8442 = _T_8440 == 1'h0; // @[LoadQueue.scala 132:9:@11905.4]
  assign storesToCheck_3_4 = _T_2318 ? _T_8435 : _T_8442; // @[LoadQueue.scala 131:10:@11906.4]
  assign _T_8448 = 4'h5 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11909.4]
  assign _T_8449 = _T_6200 & _T_8448; // @[LoadQueue.scala 131:72:@11910.4]
  assign _T_8451 = offsetQ_3 < 4'h5; // @[LoadQueue.scala 132:33:@11911.4]
  assign _T_8454 = _T_8451 & _T_6209; // @[LoadQueue.scala 132:41:@11913.4]
  assign _T_8456 = _T_8454 == 1'h0; // @[LoadQueue.scala 132:9:@11914.4]
  assign storesToCheck_3_5 = _T_2318 ? _T_8449 : _T_8456; // @[LoadQueue.scala 131:10:@11915.4]
  assign _T_8462 = 4'h6 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11918.4]
  assign _T_8463 = _T_6217 & _T_8462; // @[LoadQueue.scala 131:72:@11919.4]
  assign _T_8465 = offsetQ_3 < 4'h6; // @[LoadQueue.scala 132:33:@11920.4]
  assign _T_8468 = _T_8465 & _T_6226; // @[LoadQueue.scala 132:41:@11922.4]
  assign _T_8470 = _T_8468 == 1'h0; // @[LoadQueue.scala 132:9:@11923.4]
  assign storesToCheck_3_6 = _T_2318 ? _T_8463 : _T_8470; // @[LoadQueue.scala 131:10:@11924.4]
  assign _T_8476 = 4'h7 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11927.4]
  assign _T_8477 = _T_6234 & _T_8476; // @[LoadQueue.scala 131:72:@11928.4]
  assign _T_8479 = offsetQ_3 < 4'h7; // @[LoadQueue.scala 132:33:@11929.4]
  assign _T_8482 = _T_8479 & _T_6243; // @[LoadQueue.scala 132:41:@11931.4]
  assign _T_8484 = _T_8482 == 1'h0; // @[LoadQueue.scala 132:9:@11932.4]
  assign storesToCheck_3_7 = _T_2318 ? _T_8477 : _T_8484; // @[LoadQueue.scala 131:10:@11933.4]
  assign _T_8490 = 4'h8 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11936.4]
  assign _T_8491 = _T_6251 & _T_8490; // @[LoadQueue.scala 131:72:@11937.4]
  assign _T_8493 = offsetQ_3 < 4'h8; // @[LoadQueue.scala 132:33:@11938.4]
  assign _T_8496 = _T_8493 & _T_6260; // @[LoadQueue.scala 132:41:@11940.4]
  assign _T_8498 = _T_8496 == 1'h0; // @[LoadQueue.scala 132:9:@11941.4]
  assign storesToCheck_3_8 = _T_2318 ? _T_8491 : _T_8498; // @[LoadQueue.scala 131:10:@11942.4]
  assign _T_8504 = 4'h9 <= offsetQ_3; // @[LoadQueue.scala 131:81:@11945.4]
  assign _T_8505 = _T_6268 & _T_8504; // @[LoadQueue.scala 131:72:@11946.4]
  assign _T_8507 = offsetQ_3 < 4'h9; // @[LoadQueue.scala 132:33:@11947.4]
  assign _T_8510 = _T_8507 & _T_6277; // @[LoadQueue.scala 132:41:@11949.4]
  assign _T_8512 = _T_8510 == 1'h0; // @[LoadQueue.scala 132:9:@11950.4]
  assign storesToCheck_3_9 = _T_2318 ? _T_8505 : _T_8512; // @[LoadQueue.scala 131:10:@11951.4]
  assign _T_8518 = 4'ha <= offsetQ_3; // @[LoadQueue.scala 131:81:@11954.4]
  assign _T_8519 = _T_6285 & _T_8518; // @[LoadQueue.scala 131:72:@11955.4]
  assign _T_8521 = offsetQ_3 < 4'ha; // @[LoadQueue.scala 132:33:@11956.4]
  assign _T_8524 = _T_8521 & _T_6294; // @[LoadQueue.scala 132:41:@11958.4]
  assign _T_8526 = _T_8524 == 1'h0; // @[LoadQueue.scala 132:9:@11959.4]
  assign storesToCheck_3_10 = _T_2318 ? _T_8519 : _T_8526; // @[LoadQueue.scala 131:10:@11960.4]
  assign _T_8532 = 4'hb <= offsetQ_3; // @[LoadQueue.scala 131:81:@11963.4]
  assign _T_8533 = _T_6302 & _T_8532; // @[LoadQueue.scala 131:72:@11964.4]
  assign _T_8535 = offsetQ_3 < 4'hb; // @[LoadQueue.scala 132:33:@11965.4]
  assign _T_8538 = _T_8535 & _T_6311; // @[LoadQueue.scala 132:41:@11967.4]
  assign _T_8540 = _T_8538 == 1'h0; // @[LoadQueue.scala 132:9:@11968.4]
  assign storesToCheck_3_11 = _T_2318 ? _T_8533 : _T_8540; // @[LoadQueue.scala 131:10:@11969.4]
  assign _T_8546 = 4'hc <= offsetQ_3; // @[LoadQueue.scala 131:81:@11972.4]
  assign _T_8547 = _T_6319 & _T_8546; // @[LoadQueue.scala 131:72:@11973.4]
  assign _T_8549 = offsetQ_3 < 4'hc; // @[LoadQueue.scala 132:33:@11974.4]
  assign _T_8552 = _T_8549 & _T_6328; // @[LoadQueue.scala 132:41:@11976.4]
  assign _T_8554 = _T_8552 == 1'h0; // @[LoadQueue.scala 132:9:@11977.4]
  assign storesToCheck_3_12 = _T_2318 ? _T_8547 : _T_8554; // @[LoadQueue.scala 131:10:@11978.4]
  assign _T_8560 = 4'hd <= offsetQ_3; // @[LoadQueue.scala 131:81:@11981.4]
  assign _T_8561 = _T_6336 & _T_8560; // @[LoadQueue.scala 131:72:@11982.4]
  assign _T_8563 = offsetQ_3 < 4'hd; // @[LoadQueue.scala 132:33:@11983.4]
  assign _T_8566 = _T_8563 & _T_6345; // @[LoadQueue.scala 132:41:@11985.4]
  assign _T_8568 = _T_8566 == 1'h0; // @[LoadQueue.scala 132:9:@11986.4]
  assign storesToCheck_3_13 = _T_2318 ? _T_8561 : _T_8568; // @[LoadQueue.scala 131:10:@11987.4]
  assign _T_8574 = 4'he <= offsetQ_3; // @[LoadQueue.scala 131:81:@11990.4]
  assign _T_8575 = _T_6353 & _T_8574; // @[LoadQueue.scala 131:72:@11991.4]
  assign _T_8577 = offsetQ_3 < 4'he; // @[LoadQueue.scala 132:33:@11992.4]
  assign _T_8580 = _T_8577 & _T_6362; // @[LoadQueue.scala 132:41:@11994.4]
  assign _T_8582 = _T_8580 == 1'h0; // @[LoadQueue.scala 132:9:@11995.4]
  assign storesToCheck_3_14 = _T_2318 ? _T_8575 : _T_8582; // @[LoadQueue.scala 131:10:@11996.4]
  assign _T_8588 = 4'hf <= offsetQ_3; // @[LoadQueue.scala 131:81:@11999.4]
  assign storesToCheck_3_15 = _T_2318 ? _T_8588 : 1'h1; // @[LoadQueue.scala 131:10:@12005.4]
  assign storesToCheck_4_0 = _T_2348 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12047.4]
  assign _T_8638 = 4'h1 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12050.4]
  assign _T_8639 = _T_6132 & _T_8638; // @[LoadQueue.scala 131:72:@12051.4]
  assign _T_8641 = offsetQ_4 < 4'h1; // @[LoadQueue.scala 132:33:@12052.4]
  assign _T_8644 = _T_8641 & _T_6141; // @[LoadQueue.scala 132:41:@12054.4]
  assign _T_8646 = _T_8644 == 1'h0; // @[LoadQueue.scala 132:9:@12055.4]
  assign storesToCheck_4_1 = _T_2348 ? _T_8639 : _T_8646; // @[LoadQueue.scala 131:10:@12056.4]
  assign _T_8652 = 4'h2 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12059.4]
  assign _T_8653 = _T_6149 & _T_8652; // @[LoadQueue.scala 131:72:@12060.4]
  assign _T_8655 = offsetQ_4 < 4'h2; // @[LoadQueue.scala 132:33:@12061.4]
  assign _T_8658 = _T_8655 & _T_6158; // @[LoadQueue.scala 132:41:@12063.4]
  assign _T_8660 = _T_8658 == 1'h0; // @[LoadQueue.scala 132:9:@12064.4]
  assign storesToCheck_4_2 = _T_2348 ? _T_8653 : _T_8660; // @[LoadQueue.scala 131:10:@12065.4]
  assign _T_8666 = 4'h3 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12068.4]
  assign _T_8667 = _T_6166 & _T_8666; // @[LoadQueue.scala 131:72:@12069.4]
  assign _T_8669 = offsetQ_4 < 4'h3; // @[LoadQueue.scala 132:33:@12070.4]
  assign _T_8672 = _T_8669 & _T_6175; // @[LoadQueue.scala 132:41:@12072.4]
  assign _T_8674 = _T_8672 == 1'h0; // @[LoadQueue.scala 132:9:@12073.4]
  assign storesToCheck_4_3 = _T_2348 ? _T_8667 : _T_8674; // @[LoadQueue.scala 131:10:@12074.4]
  assign _T_8680 = 4'h4 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12077.4]
  assign _T_8681 = _T_6183 & _T_8680; // @[LoadQueue.scala 131:72:@12078.4]
  assign _T_8683 = offsetQ_4 < 4'h4; // @[LoadQueue.scala 132:33:@12079.4]
  assign _T_8686 = _T_8683 & _T_6192; // @[LoadQueue.scala 132:41:@12081.4]
  assign _T_8688 = _T_8686 == 1'h0; // @[LoadQueue.scala 132:9:@12082.4]
  assign storesToCheck_4_4 = _T_2348 ? _T_8681 : _T_8688; // @[LoadQueue.scala 131:10:@12083.4]
  assign _T_8694 = 4'h5 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12086.4]
  assign _T_8695 = _T_6200 & _T_8694; // @[LoadQueue.scala 131:72:@12087.4]
  assign _T_8697 = offsetQ_4 < 4'h5; // @[LoadQueue.scala 132:33:@12088.4]
  assign _T_8700 = _T_8697 & _T_6209; // @[LoadQueue.scala 132:41:@12090.4]
  assign _T_8702 = _T_8700 == 1'h0; // @[LoadQueue.scala 132:9:@12091.4]
  assign storesToCheck_4_5 = _T_2348 ? _T_8695 : _T_8702; // @[LoadQueue.scala 131:10:@12092.4]
  assign _T_8708 = 4'h6 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12095.4]
  assign _T_8709 = _T_6217 & _T_8708; // @[LoadQueue.scala 131:72:@12096.4]
  assign _T_8711 = offsetQ_4 < 4'h6; // @[LoadQueue.scala 132:33:@12097.4]
  assign _T_8714 = _T_8711 & _T_6226; // @[LoadQueue.scala 132:41:@12099.4]
  assign _T_8716 = _T_8714 == 1'h0; // @[LoadQueue.scala 132:9:@12100.4]
  assign storesToCheck_4_6 = _T_2348 ? _T_8709 : _T_8716; // @[LoadQueue.scala 131:10:@12101.4]
  assign _T_8722 = 4'h7 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12104.4]
  assign _T_8723 = _T_6234 & _T_8722; // @[LoadQueue.scala 131:72:@12105.4]
  assign _T_8725 = offsetQ_4 < 4'h7; // @[LoadQueue.scala 132:33:@12106.4]
  assign _T_8728 = _T_8725 & _T_6243; // @[LoadQueue.scala 132:41:@12108.4]
  assign _T_8730 = _T_8728 == 1'h0; // @[LoadQueue.scala 132:9:@12109.4]
  assign storesToCheck_4_7 = _T_2348 ? _T_8723 : _T_8730; // @[LoadQueue.scala 131:10:@12110.4]
  assign _T_8736 = 4'h8 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12113.4]
  assign _T_8737 = _T_6251 & _T_8736; // @[LoadQueue.scala 131:72:@12114.4]
  assign _T_8739 = offsetQ_4 < 4'h8; // @[LoadQueue.scala 132:33:@12115.4]
  assign _T_8742 = _T_8739 & _T_6260; // @[LoadQueue.scala 132:41:@12117.4]
  assign _T_8744 = _T_8742 == 1'h0; // @[LoadQueue.scala 132:9:@12118.4]
  assign storesToCheck_4_8 = _T_2348 ? _T_8737 : _T_8744; // @[LoadQueue.scala 131:10:@12119.4]
  assign _T_8750 = 4'h9 <= offsetQ_4; // @[LoadQueue.scala 131:81:@12122.4]
  assign _T_8751 = _T_6268 & _T_8750; // @[LoadQueue.scala 131:72:@12123.4]
  assign _T_8753 = offsetQ_4 < 4'h9; // @[LoadQueue.scala 132:33:@12124.4]
  assign _T_8756 = _T_8753 & _T_6277; // @[LoadQueue.scala 132:41:@12126.4]
  assign _T_8758 = _T_8756 == 1'h0; // @[LoadQueue.scala 132:9:@12127.4]
  assign storesToCheck_4_9 = _T_2348 ? _T_8751 : _T_8758; // @[LoadQueue.scala 131:10:@12128.4]
  assign _T_8764 = 4'ha <= offsetQ_4; // @[LoadQueue.scala 131:81:@12131.4]
  assign _T_8765 = _T_6285 & _T_8764; // @[LoadQueue.scala 131:72:@12132.4]
  assign _T_8767 = offsetQ_4 < 4'ha; // @[LoadQueue.scala 132:33:@12133.4]
  assign _T_8770 = _T_8767 & _T_6294; // @[LoadQueue.scala 132:41:@12135.4]
  assign _T_8772 = _T_8770 == 1'h0; // @[LoadQueue.scala 132:9:@12136.4]
  assign storesToCheck_4_10 = _T_2348 ? _T_8765 : _T_8772; // @[LoadQueue.scala 131:10:@12137.4]
  assign _T_8778 = 4'hb <= offsetQ_4; // @[LoadQueue.scala 131:81:@12140.4]
  assign _T_8779 = _T_6302 & _T_8778; // @[LoadQueue.scala 131:72:@12141.4]
  assign _T_8781 = offsetQ_4 < 4'hb; // @[LoadQueue.scala 132:33:@12142.4]
  assign _T_8784 = _T_8781 & _T_6311; // @[LoadQueue.scala 132:41:@12144.4]
  assign _T_8786 = _T_8784 == 1'h0; // @[LoadQueue.scala 132:9:@12145.4]
  assign storesToCheck_4_11 = _T_2348 ? _T_8779 : _T_8786; // @[LoadQueue.scala 131:10:@12146.4]
  assign _T_8792 = 4'hc <= offsetQ_4; // @[LoadQueue.scala 131:81:@12149.4]
  assign _T_8793 = _T_6319 & _T_8792; // @[LoadQueue.scala 131:72:@12150.4]
  assign _T_8795 = offsetQ_4 < 4'hc; // @[LoadQueue.scala 132:33:@12151.4]
  assign _T_8798 = _T_8795 & _T_6328; // @[LoadQueue.scala 132:41:@12153.4]
  assign _T_8800 = _T_8798 == 1'h0; // @[LoadQueue.scala 132:9:@12154.4]
  assign storesToCheck_4_12 = _T_2348 ? _T_8793 : _T_8800; // @[LoadQueue.scala 131:10:@12155.4]
  assign _T_8806 = 4'hd <= offsetQ_4; // @[LoadQueue.scala 131:81:@12158.4]
  assign _T_8807 = _T_6336 & _T_8806; // @[LoadQueue.scala 131:72:@12159.4]
  assign _T_8809 = offsetQ_4 < 4'hd; // @[LoadQueue.scala 132:33:@12160.4]
  assign _T_8812 = _T_8809 & _T_6345; // @[LoadQueue.scala 132:41:@12162.4]
  assign _T_8814 = _T_8812 == 1'h0; // @[LoadQueue.scala 132:9:@12163.4]
  assign storesToCheck_4_13 = _T_2348 ? _T_8807 : _T_8814; // @[LoadQueue.scala 131:10:@12164.4]
  assign _T_8820 = 4'he <= offsetQ_4; // @[LoadQueue.scala 131:81:@12167.4]
  assign _T_8821 = _T_6353 & _T_8820; // @[LoadQueue.scala 131:72:@12168.4]
  assign _T_8823 = offsetQ_4 < 4'he; // @[LoadQueue.scala 132:33:@12169.4]
  assign _T_8826 = _T_8823 & _T_6362; // @[LoadQueue.scala 132:41:@12171.4]
  assign _T_8828 = _T_8826 == 1'h0; // @[LoadQueue.scala 132:9:@12172.4]
  assign storesToCheck_4_14 = _T_2348 ? _T_8821 : _T_8828; // @[LoadQueue.scala 131:10:@12173.4]
  assign _T_8834 = 4'hf <= offsetQ_4; // @[LoadQueue.scala 131:81:@12176.4]
  assign storesToCheck_4_15 = _T_2348 ? _T_8834 : 1'h1; // @[LoadQueue.scala 131:10:@12182.4]
  assign storesToCheck_5_0 = _T_2378 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12224.4]
  assign _T_8884 = 4'h1 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12227.4]
  assign _T_8885 = _T_6132 & _T_8884; // @[LoadQueue.scala 131:72:@12228.4]
  assign _T_8887 = offsetQ_5 < 4'h1; // @[LoadQueue.scala 132:33:@12229.4]
  assign _T_8890 = _T_8887 & _T_6141; // @[LoadQueue.scala 132:41:@12231.4]
  assign _T_8892 = _T_8890 == 1'h0; // @[LoadQueue.scala 132:9:@12232.4]
  assign storesToCheck_5_1 = _T_2378 ? _T_8885 : _T_8892; // @[LoadQueue.scala 131:10:@12233.4]
  assign _T_8898 = 4'h2 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12236.4]
  assign _T_8899 = _T_6149 & _T_8898; // @[LoadQueue.scala 131:72:@12237.4]
  assign _T_8901 = offsetQ_5 < 4'h2; // @[LoadQueue.scala 132:33:@12238.4]
  assign _T_8904 = _T_8901 & _T_6158; // @[LoadQueue.scala 132:41:@12240.4]
  assign _T_8906 = _T_8904 == 1'h0; // @[LoadQueue.scala 132:9:@12241.4]
  assign storesToCheck_5_2 = _T_2378 ? _T_8899 : _T_8906; // @[LoadQueue.scala 131:10:@12242.4]
  assign _T_8912 = 4'h3 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12245.4]
  assign _T_8913 = _T_6166 & _T_8912; // @[LoadQueue.scala 131:72:@12246.4]
  assign _T_8915 = offsetQ_5 < 4'h3; // @[LoadQueue.scala 132:33:@12247.4]
  assign _T_8918 = _T_8915 & _T_6175; // @[LoadQueue.scala 132:41:@12249.4]
  assign _T_8920 = _T_8918 == 1'h0; // @[LoadQueue.scala 132:9:@12250.4]
  assign storesToCheck_5_3 = _T_2378 ? _T_8913 : _T_8920; // @[LoadQueue.scala 131:10:@12251.4]
  assign _T_8926 = 4'h4 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12254.4]
  assign _T_8927 = _T_6183 & _T_8926; // @[LoadQueue.scala 131:72:@12255.4]
  assign _T_8929 = offsetQ_5 < 4'h4; // @[LoadQueue.scala 132:33:@12256.4]
  assign _T_8932 = _T_8929 & _T_6192; // @[LoadQueue.scala 132:41:@12258.4]
  assign _T_8934 = _T_8932 == 1'h0; // @[LoadQueue.scala 132:9:@12259.4]
  assign storesToCheck_5_4 = _T_2378 ? _T_8927 : _T_8934; // @[LoadQueue.scala 131:10:@12260.4]
  assign _T_8940 = 4'h5 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12263.4]
  assign _T_8941 = _T_6200 & _T_8940; // @[LoadQueue.scala 131:72:@12264.4]
  assign _T_8943 = offsetQ_5 < 4'h5; // @[LoadQueue.scala 132:33:@12265.4]
  assign _T_8946 = _T_8943 & _T_6209; // @[LoadQueue.scala 132:41:@12267.4]
  assign _T_8948 = _T_8946 == 1'h0; // @[LoadQueue.scala 132:9:@12268.4]
  assign storesToCheck_5_5 = _T_2378 ? _T_8941 : _T_8948; // @[LoadQueue.scala 131:10:@12269.4]
  assign _T_8954 = 4'h6 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12272.4]
  assign _T_8955 = _T_6217 & _T_8954; // @[LoadQueue.scala 131:72:@12273.4]
  assign _T_8957 = offsetQ_5 < 4'h6; // @[LoadQueue.scala 132:33:@12274.4]
  assign _T_8960 = _T_8957 & _T_6226; // @[LoadQueue.scala 132:41:@12276.4]
  assign _T_8962 = _T_8960 == 1'h0; // @[LoadQueue.scala 132:9:@12277.4]
  assign storesToCheck_5_6 = _T_2378 ? _T_8955 : _T_8962; // @[LoadQueue.scala 131:10:@12278.4]
  assign _T_8968 = 4'h7 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12281.4]
  assign _T_8969 = _T_6234 & _T_8968; // @[LoadQueue.scala 131:72:@12282.4]
  assign _T_8971 = offsetQ_5 < 4'h7; // @[LoadQueue.scala 132:33:@12283.4]
  assign _T_8974 = _T_8971 & _T_6243; // @[LoadQueue.scala 132:41:@12285.4]
  assign _T_8976 = _T_8974 == 1'h0; // @[LoadQueue.scala 132:9:@12286.4]
  assign storesToCheck_5_7 = _T_2378 ? _T_8969 : _T_8976; // @[LoadQueue.scala 131:10:@12287.4]
  assign _T_8982 = 4'h8 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12290.4]
  assign _T_8983 = _T_6251 & _T_8982; // @[LoadQueue.scala 131:72:@12291.4]
  assign _T_8985 = offsetQ_5 < 4'h8; // @[LoadQueue.scala 132:33:@12292.4]
  assign _T_8988 = _T_8985 & _T_6260; // @[LoadQueue.scala 132:41:@12294.4]
  assign _T_8990 = _T_8988 == 1'h0; // @[LoadQueue.scala 132:9:@12295.4]
  assign storesToCheck_5_8 = _T_2378 ? _T_8983 : _T_8990; // @[LoadQueue.scala 131:10:@12296.4]
  assign _T_8996 = 4'h9 <= offsetQ_5; // @[LoadQueue.scala 131:81:@12299.4]
  assign _T_8997 = _T_6268 & _T_8996; // @[LoadQueue.scala 131:72:@12300.4]
  assign _T_8999 = offsetQ_5 < 4'h9; // @[LoadQueue.scala 132:33:@12301.4]
  assign _T_9002 = _T_8999 & _T_6277; // @[LoadQueue.scala 132:41:@12303.4]
  assign _T_9004 = _T_9002 == 1'h0; // @[LoadQueue.scala 132:9:@12304.4]
  assign storesToCheck_5_9 = _T_2378 ? _T_8997 : _T_9004; // @[LoadQueue.scala 131:10:@12305.4]
  assign _T_9010 = 4'ha <= offsetQ_5; // @[LoadQueue.scala 131:81:@12308.4]
  assign _T_9011 = _T_6285 & _T_9010; // @[LoadQueue.scala 131:72:@12309.4]
  assign _T_9013 = offsetQ_5 < 4'ha; // @[LoadQueue.scala 132:33:@12310.4]
  assign _T_9016 = _T_9013 & _T_6294; // @[LoadQueue.scala 132:41:@12312.4]
  assign _T_9018 = _T_9016 == 1'h0; // @[LoadQueue.scala 132:9:@12313.4]
  assign storesToCheck_5_10 = _T_2378 ? _T_9011 : _T_9018; // @[LoadQueue.scala 131:10:@12314.4]
  assign _T_9024 = 4'hb <= offsetQ_5; // @[LoadQueue.scala 131:81:@12317.4]
  assign _T_9025 = _T_6302 & _T_9024; // @[LoadQueue.scala 131:72:@12318.4]
  assign _T_9027 = offsetQ_5 < 4'hb; // @[LoadQueue.scala 132:33:@12319.4]
  assign _T_9030 = _T_9027 & _T_6311; // @[LoadQueue.scala 132:41:@12321.4]
  assign _T_9032 = _T_9030 == 1'h0; // @[LoadQueue.scala 132:9:@12322.4]
  assign storesToCheck_5_11 = _T_2378 ? _T_9025 : _T_9032; // @[LoadQueue.scala 131:10:@12323.4]
  assign _T_9038 = 4'hc <= offsetQ_5; // @[LoadQueue.scala 131:81:@12326.4]
  assign _T_9039 = _T_6319 & _T_9038; // @[LoadQueue.scala 131:72:@12327.4]
  assign _T_9041 = offsetQ_5 < 4'hc; // @[LoadQueue.scala 132:33:@12328.4]
  assign _T_9044 = _T_9041 & _T_6328; // @[LoadQueue.scala 132:41:@12330.4]
  assign _T_9046 = _T_9044 == 1'h0; // @[LoadQueue.scala 132:9:@12331.4]
  assign storesToCheck_5_12 = _T_2378 ? _T_9039 : _T_9046; // @[LoadQueue.scala 131:10:@12332.4]
  assign _T_9052 = 4'hd <= offsetQ_5; // @[LoadQueue.scala 131:81:@12335.4]
  assign _T_9053 = _T_6336 & _T_9052; // @[LoadQueue.scala 131:72:@12336.4]
  assign _T_9055 = offsetQ_5 < 4'hd; // @[LoadQueue.scala 132:33:@12337.4]
  assign _T_9058 = _T_9055 & _T_6345; // @[LoadQueue.scala 132:41:@12339.4]
  assign _T_9060 = _T_9058 == 1'h0; // @[LoadQueue.scala 132:9:@12340.4]
  assign storesToCheck_5_13 = _T_2378 ? _T_9053 : _T_9060; // @[LoadQueue.scala 131:10:@12341.4]
  assign _T_9066 = 4'he <= offsetQ_5; // @[LoadQueue.scala 131:81:@12344.4]
  assign _T_9067 = _T_6353 & _T_9066; // @[LoadQueue.scala 131:72:@12345.4]
  assign _T_9069 = offsetQ_5 < 4'he; // @[LoadQueue.scala 132:33:@12346.4]
  assign _T_9072 = _T_9069 & _T_6362; // @[LoadQueue.scala 132:41:@12348.4]
  assign _T_9074 = _T_9072 == 1'h0; // @[LoadQueue.scala 132:9:@12349.4]
  assign storesToCheck_5_14 = _T_2378 ? _T_9067 : _T_9074; // @[LoadQueue.scala 131:10:@12350.4]
  assign _T_9080 = 4'hf <= offsetQ_5; // @[LoadQueue.scala 131:81:@12353.4]
  assign storesToCheck_5_15 = _T_2378 ? _T_9080 : 1'h1; // @[LoadQueue.scala 131:10:@12359.4]
  assign storesToCheck_6_0 = _T_2408 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12401.4]
  assign _T_9130 = 4'h1 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12404.4]
  assign _T_9131 = _T_6132 & _T_9130; // @[LoadQueue.scala 131:72:@12405.4]
  assign _T_9133 = offsetQ_6 < 4'h1; // @[LoadQueue.scala 132:33:@12406.4]
  assign _T_9136 = _T_9133 & _T_6141; // @[LoadQueue.scala 132:41:@12408.4]
  assign _T_9138 = _T_9136 == 1'h0; // @[LoadQueue.scala 132:9:@12409.4]
  assign storesToCheck_6_1 = _T_2408 ? _T_9131 : _T_9138; // @[LoadQueue.scala 131:10:@12410.4]
  assign _T_9144 = 4'h2 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12413.4]
  assign _T_9145 = _T_6149 & _T_9144; // @[LoadQueue.scala 131:72:@12414.4]
  assign _T_9147 = offsetQ_6 < 4'h2; // @[LoadQueue.scala 132:33:@12415.4]
  assign _T_9150 = _T_9147 & _T_6158; // @[LoadQueue.scala 132:41:@12417.4]
  assign _T_9152 = _T_9150 == 1'h0; // @[LoadQueue.scala 132:9:@12418.4]
  assign storesToCheck_6_2 = _T_2408 ? _T_9145 : _T_9152; // @[LoadQueue.scala 131:10:@12419.4]
  assign _T_9158 = 4'h3 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12422.4]
  assign _T_9159 = _T_6166 & _T_9158; // @[LoadQueue.scala 131:72:@12423.4]
  assign _T_9161 = offsetQ_6 < 4'h3; // @[LoadQueue.scala 132:33:@12424.4]
  assign _T_9164 = _T_9161 & _T_6175; // @[LoadQueue.scala 132:41:@12426.4]
  assign _T_9166 = _T_9164 == 1'h0; // @[LoadQueue.scala 132:9:@12427.4]
  assign storesToCheck_6_3 = _T_2408 ? _T_9159 : _T_9166; // @[LoadQueue.scala 131:10:@12428.4]
  assign _T_9172 = 4'h4 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12431.4]
  assign _T_9173 = _T_6183 & _T_9172; // @[LoadQueue.scala 131:72:@12432.4]
  assign _T_9175 = offsetQ_6 < 4'h4; // @[LoadQueue.scala 132:33:@12433.4]
  assign _T_9178 = _T_9175 & _T_6192; // @[LoadQueue.scala 132:41:@12435.4]
  assign _T_9180 = _T_9178 == 1'h0; // @[LoadQueue.scala 132:9:@12436.4]
  assign storesToCheck_6_4 = _T_2408 ? _T_9173 : _T_9180; // @[LoadQueue.scala 131:10:@12437.4]
  assign _T_9186 = 4'h5 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12440.4]
  assign _T_9187 = _T_6200 & _T_9186; // @[LoadQueue.scala 131:72:@12441.4]
  assign _T_9189 = offsetQ_6 < 4'h5; // @[LoadQueue.scala 132:33:@12442.4]
  assign _T_9192 = _T_9189 & _T_6209; // @[LoadQueue.scala 132:41:@12444.4]
  assign _T_9194 = _T_9192 == 1'h0; // @[LoadQueue.scala 132:9:@12445.4]
  assign storesToCheck_6_5 = _T_2408 ? _T_9187 : _T_9194; // @[LoadQueue.scala 131:10:@12446.4]
  assign _T_9200 = 4'h6 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12449.4]
  assign _T_9201 = _T_6217 & _T_9200; // @[LoadQueue.scala 131:72:@12450.4]
  assign _T_9203 = offsetQ_6 < 4'h6; // @[LoadQueue.scala 132:33:@12451.4]
  assign _T_9206 = _T_9203 & _T_6226; // @[LoadQueue.scala 132:41:@12453.4]
  assign _T_9208 = _T_9206 == 1'h0; // @[LoadQueue.scala 132:9:@12454.4]
  assign storesToCheck_6_6 = _T_2408 ? _T_9201 : _T_9208; // @[LoadQueue.scala 131:10:@12455.4]
  assign _T_9214 = 4'h7 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12458.4]
  assign _T_9215 = _T_6234 & _T_9214; // @[LoadQueue.scala 131:72:@12459.4]
  assign _T_9217 = offsetQ_6 < 4'h7; // @[LoadQueue.scala 132:33:@12460.4]
  assign _T_9220 = _T_9217 & _T_6243; // @[LoadQueue.scala 132:41:@12462.4]
  assign _T_9222 = _T_9220 == 1'h0; // @[LoadQueue.scala 132:9:@12463.4]
  assign storesToCheck_6_7 = _T_2408 ? _T_9215 : _T_9222; // @[LoadQueue.scala 131:10:@12464.4]
  assign _T_9228 = 4'h8 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12467.4]
  assign _T_9229 = _T_6251 & _T_9228; // @[LoadQueue.scala 131:72:@12468.4]
  assign _T_9231 = offsetQ_6 < 4'h8; // @[LoadQueue.scala 132:33:@12469.4]
  assign _T_9234 = _T_9231 & _T_6260; // @[LoadQueue.scala 132:41:@12471.4]
  assign _T_9236 = _T_9234 == 1'h0; // @[LoadQueue.scala 132:9:@12472.4]
  assign storesToCheck_6_8 = _T_2408 ? _T_9229 : _T_9236; // @[LoadQueue.scala 131:10:@12473.4]
  assign _T_9242 = 4'h9 <= offsetQ_6; // @[LoadQueue.scala 131:81:@12476.4]
  assign _T_9243 = _T_6268 & _T_9242; // @[LoadQueue.scala 131:72:@12477.4]
  assign _T_9245 = offsetQ_6 < 4'h9; // @[LoadQueue.scala 132:33:@12478.4]
  assign _T_9248 = _T_9245 & _T_6277; // @[LoadQueue.scala 132:41:@12480.4]
  assign _T_9250 = _T_9248 == 1'h0; // @[LoadQueue.scala 132:9:@12481.4]
  assign storesToCheck_6_9 = _T_2408 ? _T_9243 : _T_9250; // @[LoadQueue.scala 131:10:@12482.4]
  assign _T_9256 = 4'ha <= offsetQ_6; // @[LoadQueue.scala 131:81:@12485.4]
  assign _T_9257 = _T_6285 & _T_9256; // @[LoadQueue.scala 131:72:@12486.4]
  assign _T_9259 = offsetQ_6 < 4'ha; // @[LoadQueue.scala 132:33:@12487.4]
  assign _T_9262 = _T_9259 & _T_6294; // @[LoadQueue.scala 132:41:@12489.4]
  assign _T_9264 = _T_9262 == 1'h0; // @[LoadQueue.scala 132:9:@12490.4]
  assign storesToCheck_6_10 = _T_2408 ? _T_9257 : _T_9264; // @[LoadQueue.scala 131:10:@12491.4]
  assign _T_9270 = 4'hb <= offsetQ_6; // @[LoadQueue.scala 131:81:@12494.4]
  assign _T_9271 = _T_6302 & _T_9270; // @[LoadQueue.scala 131:72:@12495.4]
  assign _T_9273 = offsetQ_6 < 4'hb; // @[LoadQueue.scala 132:33:@12496.4]
  assign _T_9276 = _T_9273 & _T_6311; // @[LoadQueue.scala 132:41:@12498.4]
  assign _T_9278 = _T_9276 == 1'h0; // @[LoadQueue.scala 132:9:@12499.4]
  assign storesToCheck_6_11 = _T_2408 ? _T_9271 : _T_9278; // @[LoadQueue.scala 131:10:@12500.4]
  assign _T_9284 = 4'hc <= offsetQ_6; // @[LoadQueue.scala 131:81:@12503.4]
  assign _T_9285 = _T_6319 & _T_9284; // @[LoadQueue.scala 131:72:@12504.4]
  assign _T_9287 = offsetQ_6 < 4'hc; // @[LoadQueue.scala 132:33:@12505.4]
  assign _T_9290 = _T_9287 & _T_6328; // @[LoadQueue.scala 132:41:@12507.4]
  assign _T_9292 = _T_9290 == 1'h0; // @[LoadQueue.scala 132:9:@12508.4]
  assign storesToCheck_6_12 = _T_2408 ? _T_9285 : _T_9292; // @[LoadQueue.scala 131:10:@12509.4]
  assign _T_9298 = 4'hd <= offsetQ_6; // @[LoadQueue.scala 131:81:@12512.4]
  assign _T_9299 = _T_6336 & _T_9298; // @[LoadQueue.scala 131:72:@12513.4]
  assign _T_9301 = offsetQ_6 < 4'hd; // @[LoadQueue.scala 132:33:@12514.4]
  assign _T_9304 = _T_9301 & _T_6345; // @[LoadQueue.scala 132:41:@12516.4]
  assign _T_9306 = _T_9304 == 1'h0; // @[LoadQueue.scala 132:9:@12517.4]
  assign storesToCheck_6_13 = _T_2408 ? _T_9299 : _T_9306; // @[LoadQueue.scala 131:10:@12518.4]
  assign _T_9312 = 4'he <= offsetQ_6; // @[LoadQueue.scala 131:81:@12521.4]
  assign _T_9313 = _T_6353 & _T_9312; // @[LoadQueue.scala 131:72:@12522.4]
  assign _T_9315 = offsetQ_6 < 4'he; // @[LoadQueue.scala 132:33:@12523.4]
  assign _T_9318 = _T_9315 & _T_6362; // @[LoadQueue.scala 132:41:@12525.4]
  assign _T_9320 = _T_9318 == 1'h0; // @[LoadQueue.scala 132:9:@12526.4]
  assign storesToCheck_6_14 = _T_2408 ? _T_9313 : _T_9320; // @[LoadQueue.scala 131:10:@12527.4]
  assign _T_9326 = 4'hf <= offsetQ_6; // @[LoadQueue.scala 131:81:@12530.4]
  assign storesToCheck_6_15 = _T_2408 ? _T_9326 : 1'h1; // @[LoadQueue.scala 131:10:@12536.4]
  assign storesToCheck_7_0 = _T_2438 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12578.4]
  assign _T_9376 = 4'h1 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12581.4]
  assign _T_9377 = _T_6132 & _T_9376; // @[LoadQueue.scala 131:72:@12582.4]
  assign _T_9379 = offsetQ_7 < 4'h1; // @[LoadQueue.scala 132:33:@12583.4]
  assign _T_9382 = _T_9379 & _T_6141; // @[LoadQueue.scala 132:41:@12585.4]
  assign _T_9384 = _T_9382 == 1'h0; // @[LoadQueue.scala 132:9:@12586.4]
  assign storesToCheck_7_1 = _T_2438 ? _T_9377 : _T_9384; // @[LoadQueue.scala 131:10:@12587.4]
  assign _T_9390 = 4'h2 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12590.4]
  assign _T_9391 = _T_6149 & _T_9390; // @[LoadQueue.scala 131:72:@12591.4]
  assign _T_9393 = offsetQ_7 < 4'h2; // @[LoadQueue.scala 132:33:@12592.4]
  assign _T_9396 = _T_9393 & _T_6158; // @[LoadQueue.scala 132:41:@12594.4]
  assign _T_9398 = _T_9396 == 1'h0; // @[LoadQueue.scala 132:9:@12595.4]
  assign storesToCheck_7_2 = _T_2438 ? _T_9391 : _T_9398; // @[LoadQueue.scala 131:10:@12596.4]
  assign _T_9404 = 4'h3 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12599.4]
  assign _T_9405 = _T_6166 & _T_9404; // @[LoadQueue.scala 131:72:@12600.4]
  assign _T_9407 = offsetQ_7 < 4'h3; // @[LoadQueue.scala 132:33:@12601.4]
  assign _T_9410 = _T_9407 & _T_6175; // @[LoadQueue.scala 132:41:@12603.4]
  assign _T_9412 = _T_9410 == 1'h0; // @[LoadQueue.scala 132:9:@12604.4]
  assign storesToCheck_7_3 = _T_2438 ? _T_9405 : _T_9412; // @[LoadQueue.scala 131:10:@12605.4]
  assign _T_9418 = 4'h4 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12608.4]
  assign _T_9419 = _T_6183 & _T_9418; // @[LoadQueue.scala 131:72:@12609.4]
  assign _T_9421 = offsetQ_7 < 4'h4; // @[LoadQueue.scala 132:33:@12610.4]
  assign _T_9424 = _T_9421 & _T_6192; // @[LoadQueue.scala 132:41:@12612.4]
  assign _T_9426 = _T_9424 == 1'h0; // @[LoadQueue.scala 132:9:@12613.4]
  assign storesToCheck_7_4 = _T_2438 ? _T_9419 : _T_9426; // @[LoadQueue.scala 131:10:@12614.4]
  assign _T_9432 = 4'h5 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12617.4]
  assign _T_9433 = _T_6200 & _T_9432; // @[LoadQueue.scala 131:72:@12618.4]
  assign _T_9435 = offsetQ_7 < 4'h5; // @[LoadQueue.scala 132:33:@12619.4]
  assign _T_9438 = _T_9435 & _T_6209; // @[LoadQueue.scala 132:41:@12621.4]
  assign _T_9440 = _T_9438 == 1'h0; // @[LoadQueue.scala 132:9:@12622.4]
  assign storesToCheck_7_5 = _T_2438 ? _T_9433 : _T_9440; // @[LoadQueue.scala 131:10:@12623.4]
  assign _T_9446 = 4'h6 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12626.4]
  assign _T_9447 = _T_6217 & _T_9446; // @[LoadQueue.scala 131:72:@12627.4]
  assign _T_9449 = offsetQ_7 < 4'h6; // @[LoadQueue.scala 132:33:@12628.4]
  assign _T_9452 = _T_9449 & _T_6226; // @[LoadQueue.scala 132:41:@12630.4]
  assign _T_9454 = _T_9452 == 1'h0; // @[LoadQueue.scala 132:9:@12631.4]
  assign storesToCheck_7_6 = _T_2438 ? _T_9447 : _T_9454; // @[LoadQueue.scala 131:10:@12632.4]
  assign _T_9460 = 4'h7 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12635.4]
  assign _T_9461 = _T_6234 & _T_9460; // @[LoadQueue.scala 131:72:@12636.4]
  assign _T_9463 = offsetQ_7 < 4'h7; // @[LoadQueue.scala 132:33:@12637.4]
  assign _T_9466 = _T_9463 & _T_6243; // @[LoadQueue.scala 132:41:@12639.4]
  assign _T_9468 = _T_9466 == 1'h0; // @[LoadQueue.scala 132:9:@12640.4]
  assign storesToCheck_7_7 = _T_2438 ? _T_9461 : _T_9468; // @[LoadQueue.scala 131:10:@12641.4]
  assign _T_9474 = 4'h8 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12644.4]
  assign _T_9475 = _T_6251 & _T_9474; // @[LoadQueue.scala 131:72:@12645.4]
  assign _T_9477 = offsetQ_7 < 4'h8; // @[LoadQueue.scala 132:33:@12646.4]
  assign _T_9480 = _T_9477 & _T_6260; // @[LoadQueue.scala 132:41:@12648.4]
  assign _T_9482 = _T_9480 == 1'h0; // @[LoadQueue.scala 132:9:@12649.4]
  assign storesToCheck_7_8 = _T_2438 ? _T_9475 : _T_9482; // @[LoadQueue.scala 131:10:@12650.4]
  assign _T_9488 = 4'h9 <= offsetQ_7; // @[LoadQueue.scala 131:81:@12653.4]
  assign _T_9489 = _T_6268 & _T_9488; // @[LoadQueue.scala 131:72:@12654.4]
  assign _T_9491 = offsetQ_7 < 4'h9; // @[LoadQueue.scala 132:33:@12655.4]
  assign _T_9494 = _T_9491 & _T_6277; // @[LoadQueue.scala 132:41:@12657.4]
  assign _T_9496 = _T_9494 == 1'h0; // @[LoadQueue.scala 132:9:@12658.4]
  assign storesToCheck_7_9 = _T_2438 ? _T_9489 : _T_9496; // @[LoadQueue.scala 131:10:@12659.4]
  assign _T_9502 = 4'ha <= offsetQ_7; // @[LoadQueue.scala 131:81:@12662.4]
  assign _T_9503 = _T_6285 & _T_9502; // @[LoadQueue.scala 131:72:@12663.4]
  assign _T_9505 = offsetQ_7 < 4'ha; // @[LoadQueue.scala 132:33:@12664.4]
  assign _T_9508 = _T_9505 & _T_6294; // @[LoadQueue.scala 132:41:@12666.4]
  assign _T_9510 = _T_9508 == 1'h0; // @[LoadQueue.scala 132:9:@12667.4]
  assign storesToCheck_7_10 = _T_2438 ? _T_9503 : _T_9510; // @[LoadQueue.scala 131:10:@12668.4]
  assign _T_9516 = 4'hb <= offsetQ_7; // @[LoadQueue.scala 131:81:@12671.4]
  assign _T_9517 = _T_6302 & _T_9516; // @[LoadQueue.scala 131:72:@12672.4]
  assign _T_9519 = offsetQ_7 < 4'hb; // @[LoadQueue.scala 132:33:@12673.4]
  assign _T_9522 = _T_9519 & _T_6311; // @[LoadQueue.scala 132:41:@12675.4]
  assign _T_9524 = _T_9522 == 1'h0; // @[LoadQueue.scala 132:9:@12676.4]
  assign storesToCheck_7_11 = _T_2438 ? _T_9517 : _T_9524; // @[LoadQueue.scala 131:10:@12677.4]
  assign _T_9530 = 4'hc <= offsetQ_7; // @[LoadQueue.scala 131:81:@12680.4]
  assign _T_9531 = _T_6319 & _T_9530; // @[LoadQueue.scala 131:72:@12681.4]
  assign _T_9533 = offsetQ_7 < 4'hc; // @[LoadQueue.scala 132:33:@12682.4]
  assign _T_9536 = _T_9533 & _T_6328; // @[LoadQueue.scala 132:41:@12684.4]
  assign _T_9538 = _T_9536 == 1'h0; // @[LoadQueue.scala 132:9:@12685.4]
  assign storesToCheck_7_12 = _T_2438 ? _T_9531 : _T_9538; // @[LoadQueue.scala 131:10:@12686.4]
  assign _T_9544 = 4'hd <= offsetQ_7; // @[LoadQueue.scala 131:81:@12689.4]
  assign _T_9545 = _T_6336 & _T_9544; // @[LoadQueue.scala 131:72:@12690.4]
  assign _T_9547 = offsetQ_7 < 4'hd; // @[LoadQueue.scala 132:33:@12691.4]
  assign _T_9550 = _T_9547 & _T_6345; // @[LoadQueue.scala 132:41:@12693.4]
  assign _T_9552 = _T_9550 == 1'h0; // @[LoadQueue.scala 132:9:@12694.4]
  assign storesToCheck_7_13 = _T_2438 ? _T_9545 : _T_9552; // @[LoadQueue.scala 131:10:@12695.4]
  assign _T_9558 = 4'he <= offsetQ_7; // @[LoadQueue.scala 131:81:@12698.4]
  assign _T_9559 = _T_6353 & _T_9558; // @[LoadQueue.scala 131:72:@12699.4]
  assign _T_9561 = offsetQ_7 < 4'he; // @[LoadQueue.scala 132:33:@12700.4]
  assign _T_9564 = _T_9561 & _T_6362; // @[LoadQueue.scala 132:41:@12702.4]
  assign _T_9566 = _T_9564 == 1'h0; // @[LoadQueue.scala 132:9:@12703.4]
  assign storesToCheck_7_14 = _T_2438 ? _T_9559 : _T_9566; // @[LoadQueue.scala 131:10:@12704.4]
  assign _T_9572 = 4'hf <= offsetQ_7; // @[LoadQueue.scala 131:81:@12707.4]
  assign storesToCheck_7_15 = _T_2438 ? _T_9572 : 1'h1; // @[LoadQueue.scala 131:10:@12713.4]
  assign storesToCheck_8_0 = _T_2468 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12755.4]
  assign _T_9622 = 4'h1 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12758.4]
  assign _T_9623 = _T_6132 & _T_9622; // @[LoadQueue.scala 131:72:@12759.4]
  assign _T_9625 = offsetQ_8 < 4'h1; // @[LoadQueue.scala 132:33:@12760.4]
  assign _T_9628 = _T_9625 & _T_6141; // @[LoadQueue.scala 132:41:@12762.4]
  assign _T_9630 = _T_9628 == 1'h0; // @[LoadQueue.scala 132:9:@12763.4]
  assign storesToCheck_8_1 = _T_2468 ? _T_9623 : _T_9630; // @[LoadQueue.scala 131:10:@12764.4]
  assign _T_9636 = 4'h2 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12767.4]
  assign _T_9637 = _T_6149 & _T_9636; // @[LoadQueue.scala 131:72:@12768.4]
  assign _T_9639 = offsetQ_8 < 4'h2; // @[LoadQueue.scala 132:33:@12769.4]
  assign _T_9642 = _T_9639 & _T_6158; // @[LoadQueue.scala 132:41:@12771.4]
  assign _T_9644 = _T_9642 == 1'h0; // @[LoadQueue.scala 132:9:@12772.4]
  assign storesToCheck_8_2 = _T_2468 ? _T_9637 : _T_9644; // @[LoadQueue.scala 131:10:@12773.4]
  assign _T_9650 = 4'h3 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12776.4]
  assign _T_9651 = _T_6166 & _T_9650; // @[LoadQueue.scala 131:72:@12777.4]
  assign _T_9653 = offsetQ_8 < 4'h3; // @[LoadQueue.scala 132:33:@12778.4]
  assign _T_9656 = _T_9653 & _T_6175; // @[LoadQueue.scala 132:41:@12780.4]
  assign _T_9658 = _T_9656 == 1'h0; // @[LoadQueue.scala 132:9:@12781.4]
  assign storesToCheck_8_3 = _T_2468 ? _T_9651 : _T_9658; // @[LoadQueue.scala 131:10:@12782.4]
  assign _T_9664 = 4'h4 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12785.4]
  assign _T_9665 = _T_6183 & _T_9664; // @[LoadQueue.scala 131:72:@12786.4]
  assign _T_9667 = offsetQ_8 < 4'h4; // @[LoadQueue.scala 132:33:@12787.4]
  assign _T_9670 = _T_9667 & _T_6192; // @[LoadQueue.scala 132:41:@12789.4]
  assign _T_9672 = _T_9670 == 1'h0; // @[LoadQueue.scala 132:9:@12790.4]
  assign storesToCheck_8_4 = _T_2468 ? _T_9665 : _T_9672; // @[LoadQueue.scala 131:10:@12791.4]
  assign _T_9678 = 4'h5 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12794.4]
  assign _T_9679 = _T_6200 & _T_9678; // @[LoadQueue.scala 131:72:@12795.4]
  assign _T_9681 = offsetQ_8 < 4'h5; // @[LoadQueue.scala 132:33:@12796.4]
  assign _T_9684 = _T_9681 & _T_6209; // @[LoadQueue.scala 132:41:@12798.4]
  assign _T_9686 = _T_9684 == 1'h0; // @[LoadQueue.scala 132:9:@12799.4]
  assign storesToCheck_8_5 = _T_2468 ? _T_9679 : _T_9686; // @[LoadQueue.scala 131:10:@12800.4]
  assign _T_9692 = 4'h6 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12803.4]
  assign _T_9693 = _T_6217 & _T_9692; // @[LoadQueue.scala 131:72:@12804.4]
  assign _T_9695 = offsetQ_8 < 4'h6; // @[LoadQueue.scala 132:33:@12805.4]
  assign _T_9698 = _T_9695 & _T_6226; // @[LoadQueue.scala 132:41:@12807.4]
  assign _T_9700 = _T_9698 == 1'h0; // @[LoadQueue.scala 132:9:@12808.4]
  assign storesToCheck_8_6 = _T_2468 ? _T_9693 : _T_9700; // @[LoadQueue.scala 131:10:@12809.4]
  assign _T_9706 = 4'h7 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12812.4]
  assign _T_9707 = _T_6234 & _T_9706; // @[LoadQueue.scala 131:72:@12813.4]
  assign _T_9709 = offsetQ_8 < 4'h7; // @[LoadQueue.scala 132:33:@12814.4]
  assign _T_9712 = _T_9709 & _T_6243; // @[LoadQueue.scala 132:41:@12816.4]
  assign _T_9714 = _T_9712 == 1'h0; // @[LoadQueue.scala 132:9:@12817.4]
  assign storesToCheck_8_7 = _T_2468 ? _T_9707 : _T_9714; // @[LoadQueue.scala 131:10:@12818.4]
  assign _T_9720 = 4'h8 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12821.4]
  assign _T_9721 = _T_6251 & _T_9720; // @[LoadQueue.scala 131:72:@12822.4]
  assign _T_9723 = offsetQ_8 < 4'h8; // @[LoadQueue.scala 132:33:@12823.4]
  assign _T_9726 = _T_9723 & _T_6260; // @[LoadQueue.scala 132:41:@12825.4]
  assign _T_9728 = _T_9726 == 1'h0; // @[LoadQueue.scala 132:9:@12826.4]
  assign storesToCheck_8_8 = _T_2468 ? _T_9721 : _T_9728; // @[LoadQueue.scala 131:10:@12827.4]
  assign _T_9734 = 4'h9 <= offsetQ_8; // @[LoadQueue.scala 131:81:@12830.4]
  assign _T_9735 = _T_6268 & _T_9734; // @[LoadQueue.scala 131:72:@12831.4]
  assign _T_9737 = offsetQ_8 < 4'h9; // @[LoadQueue.scala 132:33:@12832.4]
  assign _T_9740 = _T_9737 & _T_6277; // @[LoadQueue.scala 132:41:@12834.4]
  assign _T_9742 = _T_9740 == 1'h0; // @[LoadQueue.scala 132:9:@12835.4]
  assign storesToCheck_8_9 = _T_2468 ? _T_9735 : _T_9742; // @[LoadQueue.scala 131:10:@12836.4]
  assign _T_9748 = 4'ha <= offsetQ_8; // @[LoadQueue.scala 131:81:@12839.4]
  assign _T_9749 = _T_6285 & _T_9748; // @[LoadQueue.scala 131:72:@12840.4]
  assign _T_9751 = offsetQ_8 < 4'ha; // @[LoadQueue.scala 132:33:@12841.4]
  assign _T_9754 = _T_9751 & _T_6294; // @[LoadQueue.scala 132:41:@12843.4]
  assign _T_9756 = _T_9754 == 1'h0; // @[LoadQueue.scala 132:9:@12844.4]
  assign storesToCheck_8_10 = _T_2468 ? _T_9749 : _T_9756; // @[LoadQueue.scala 131:10:@12845.4]
  assign _T_9762 = 4'hb <= offsetQ_8; // @[LoadQueue.scala 131:81:@12848.4]
  assign _T_9763 = _T_6302 & _T_9762; // @[LoadQueue.scala 131:72:@12849.4]
  assign _T_9765 = offsetQ_8 < 4'hb; // @[LoadQueue.scala 132:33:@12850.4]
  assign _T_9768 = _T_9765 & _T_6311; // @[LoadQueue.scala 132:41:@12852.4]
  assign _T_9770 = _T_9768 == 1'h0; // @[LoadQueue.scala 132:9:@12853.4]
  assign storesToCheck_8_11 = _T_2468 ? _T_9763 : _T_9770; // @[LoadQueue.scala 131:10:@12854.4]
  assign _T_9776 = 4'hc <= offsetQ_8; // @[LoadQueue.scala 131:81:@12857.4]
  assign _T_9777 = _T_6319 & _T_9776; // @[LoadQueue.scala 131:72:@12858.4]
  assign _T_9779 = offsetQ_8 < 4'hc; // @[LoadQueue.scala 132:33:@12859.4]
  assign _T_9782 = _T_9779 & _T_6328; // @[LoadQueue.scala 132:41:@12861.4]
  assign _T_9784 = _T_9782 == 1'h0; // @[LoadQueue.scala 132:9:@12862.4]
  assign storesToCheck_8_12 = _T_2468 ? _T_9777 : _T_9784; // @[LoadQueue.scala 131:10:@12863.4]
  assign _T_9790 = 4'hd <= offsetQ_8; // @[LoadQueue.scala 131:81:@12866.4]
  assign _T_9791 = _T_6336 & _T_9790; // @[LoadQueue.scala 131:72:@12867.4]
  assign _T_9793 = offsetQ_8 < 4'hd; // @[LoadQueue.scala 132:33:@12868.4]
  assign _T_9796 = _T_9793 & _T_6345; // @[LoadQueue.scala 132:41:@12870.4]
  assign _T_9798 = _T_9796 == 1'h0; // @[LoadQueue.scala 132:9:@12871.4]
  assign storesToCheck_8_13 = _T_2468 ? _T_9791 : _T_9798; // @[LoadQueue.scala 131:10:@12872.4]
  assign _T_9804 = 4'he <= offsetQ_8; // @[LoadQueue.scala 131:81:@12875.4]
  assign _T_9805 = _T_6353 & _T_9804; // @[LoadQueue.scala 131:72:@12876.4]
  assign _T_9807 = offsetQ_8 < 4'he; // @[LoadQueue.scala 132:33:@12877.4]
  assign _T_9810 = _T_9807 & _T_6362; // @[LoadQueue.scala 132:41:@12879.4]
  assign _T_9812 = _T_9810 == 1'h0; // @[LoadQueue.scala 132:9:@12880.4]
  assign storesToCheck_8_14 = _T_2468 ? _T_9805 : _T_9812; // @[LoadQueue.scala 131:10:@12881.4]
  assign _T_9818 = 4'hf <= offsetQ_8; // @[LoadQueue.scala 131:81:@12884.4]
  assign storesToCheck_8_15 = _T_2468 ? _T_9818 : 1'h1; // @[LoadQueue.scala 131:10:@12890.4]
  assign storesToCheck_9_0 = _T_2498 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@12932.4]
  assign _T_9868 = 4'h1 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12935.4]
  assign _T_9869 = _T_6132 & _T_9868; // @[LoadQueue.scala 131:72:@12936.4]
  assign _T_9871 = offsetQ_9 < 4'h1; // @[LoadQueue.scala 132:33:@12937.4]
  assign _T_9874 = _T_9871 & _T_6141; // @[LoadQueue.scala 132:41:@12939.4]
  assign _T_9876 = _T_9874 == 1'h0; // @[LoadQueue.scala 132:9:@12940.4]
  assign storesToCheck_9_1 = _T_2498 ? _T_9869 : _T_9876; // @[LoadQueue.scala 131:10:@12941.4]
  assign _T_9882 = 4'h2 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12944.4]
  assign _T_9883 = _T_6149 & _T_9882; // @[LoadQueue.scala 131:72:@12945.4]
  assign _T_9885 = offsetQ_9 < 4'h2; // @[LoadQueue.scala 132:33:@12946.4]
  assign _T_9888 = _T_9885 & _T_6158; // @[LoadQueue.scala 132:41:@12948.4]
  assign _T_9890 = _T_9888 == 1'h0; // @[LoadQueue.scala 132:9:@12949.4]
  assign storesToCheck_9_2 = _T_2498 ? _T_9883 : _T_9890; // @[LoadQueue.scala 131:10:@12950.4]
  assign _T_9896 = 4'h3 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12953.4]
  assign _T_9897 = _T_6166 & _T_9896; // @[LoadQueue.scala 131:72:@12954.4]
  assign _T_9899 = offsetQ_9 < 4'h3; // @[LoadQueue.scala 132:33:@12955.4]
  assign _T_9902 = _T_9899 & _T_6175; // @[LoadQueue.scala 132:41:@12957.4]
  assign _T_9904 = _T_9902 == 1'h0; // @[LoadQueue.scala 132:9:@12958.4]
  assign storesToCheck_9_3 = _T_2498 ? _T_9897 : _T_9904; // @[LoadQueue.scala 131:10:@12959.4]
  assign _T_9910 = 4'h4 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12962.4]
  assign _T_9911 = _T_6183 & _T_9910; // @[LoadQueue.scala 131:72:@12963.4]
  assign _T_9913 = offsetQ_9 < 4'h4; // @[LoadQueue.scala 132:33:@12964.4]
  assign _T_9916 = _T_9913 & _T_6192; // @[LoadQueue.scala 132:41:@12966.4]
  assign _T_9918 = _T_9916 == 1'h0; // @[LoadQueue.scala 132:9:@12967.4]
  assign storesToCheck_9_4 = _T_2498 ? _T_9911 : _T_9918; // @[LoadQueue.scala 131:10:@12968.4]
  assign _T_9924 = 4'h5 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12971.4]
  assign _T_9925 = _T_6200 & _T_9924; // @[LoadQueue.scala 131:72:@12972.4]
  assign _T_9927 = offsetQ_9 < 4'h5; // @[LoadQueue.scala 132:33:@12973.4]
  assign _T_9930 = _T_9927 & _T_6209; // @[LoadQueue.scala 132:41:@12975.4]
  assign _T_9932 = _T_9930 == 1'h0; // @[LoadQueue.scala 132:9:@12976.4]
  assign storesToCheck_9_5 = _T_2498 ? _T_9925 : _T_9932; // @[LoadQueue.scala 131:10:@12977.4]
  assign _T_9938 = 4'h6 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12980.4]
  assign _T_9939 = _T_6217 & _T_9938; // @[LoadQueue.scala 131:72:@12981.4]
  assign _T_9941 = offsetQ_9 < 4'h6; // @[LoadQueue.scala 132:33:@12982.4]
  assign _T_9944 = _T_9941 & _T_6226; // @[LoadQueue.scala 132:41:@12984.4]
  assign _T_9946 = _T_9944 == 1'h0; // @[LoadQueue.scala 132:9:@12985.4]
  assign storesToCheck_9_6 = _T_2498 ? _T_9939 : _T_9946; // @[LoadQueue.scala 131:10:@12986.4]
  assign _T_9952 = 4'h7 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12989.4]
  assign _T_9953 = _T_6234 & _T_9952; // @[LoadQueue.scala 131:72:@12990.4]
  assign _T_9955 = offsetQ_9 < 4'h7; // @[LoadQueue.scala 132:33:@12991.4]
  assign _T_9958 = _T_9955 & _T_6243; // @[LoadQueue.scala 132:41:@12993.4]
  assign _T_9960 = _T_9958 == 1'h0; // @[LoadQueue.scala 132:9:@12994.4]
  assign storesToCheck_9_7 = _T_2498 ? _T_9953 : _T_9960; // @[LoadQueue.scala 131:10:@12995.4]
  assign _T_9966 = 4'h8 <= offsetQ_9; // @[LoadQueue.scala 131:81:@12998.4]
  assign _T_9967 = _T_6251 & _T_9966; // @[LoadQueue.scala 131:72:@12999.4]
  assign _T_9969 = offsetQ_9 < 4'h8; // @[LoadQueue.scala 132:33:@13000.4]
  assign _T_9972 = _T_9969 & _T_6260; // @[LoadQueue.scala 132:41:@13002.4]
  assign _T_9974 = _T_9972 == 1'h0; // @[LoadQueue.scala 132:9:@13003.4]
  assign storesToCheck_9_8 = _T_2498 ? _T_9967 : _T_9974; // @[LoadQueue.scala 131:10:@13004.4]
  assign _T_9980 = 4'h9 <= offsetQ_9; // @[LoadQueue.scala 131:81:@13007.4]
  assign _T_9981 = _T_6268 & _T_9980; // @[LoadQueue.scala 131:72:@13008.4]
  assign _T_9983 = offsetQ_9 < 4'h9; // @[LoadQueue.scala 132:33:@13009.4]
  assign _T_9986 = _T_9983 & _T_6277; // @[LoadQueue.scala 132:41:@13011.4]
  assign _T_9988 = _T_9986 == 1'h0; // @[LoadQueue.scala 132:9:@13012.4]
  assign storesToCheck_9_9 = _T_2498 ? _T_9981 : _T_9988; // @[LoadQueue.scala 131:10:@13013.4]
  assign _T_9994 = 4'ha <= offsetQ_9; // @[LoadQueue.scala 131:81:@13016.4]
  assign _T_9995 = _T_6285 & _T_9994; // @[LoadQueue.scala 131:72:@13017.4]
  assign _T_9997 = offsetQ_9 < 4'ha; // @[LoadQueue.scala 132:33:@13018.4]
  assign _T_10000 = _T_9997 & _T_6294; // @[LoadQueue.scala 132:41:@13020.4]
  assign _T_10002 = _T_10000 == 1'h0; // @[LoadQueue.scala 132:9:@13021.4]
  assign storesToCheck_9_10 = _T_2498 ? _T_9995 : _T_10002; // @[LoadQueue.scala 131:10:@13022.4]
  assign _T_10008 = 4'hb <= offsetQ_9; // @[LoadQueue.scala 131:81:@13025.4]
  assign _T_10009 = _T_6302 & _T_10008; // @[LoadQueue.scala 131:72:@13026.4]
  assign _T_10011 = offsetQ_9 < 4'hb; // @[LoadQueue.scala 132:33:@13027.4]
  assign _T_10014 = _T_10011 & _T_6311; // @[LoadQueue.scala 132:41:@13029.4]
  assign _T_10016 = _T_10014 == 1'h0; // @[LoadQueue.scala 132:9:@13030.4]
  assign storesToCheck_9_11 = _T_2498 ? _T_10009 : _T_10016; // @[LoadQueue.scala 131:10:@13031.4]
  assign _T_10022 = 4'hc <= offsetQ_9; // @[LoadQueue.scala 131:81:@13034.4]
  assign _T_10023 = _T_6319 & _T_10022; // @[LoadQueue.scala 131:72:@13035.4]
  assign _T_10025 = offsetQ_9 < 4'hc; // @[LoadQueue.scala 132:33:@13036.4]
  assign _T_10028 = _T_10025 & _T_6328; // @[LoadQueue.scala 132:41:@13038.4]
  assign _T_10030 = _T_10028 == 1'h0; // @[LoadQueue.scala 132:9:@13039.4]
  assign storesToCheck_9_12 = _T_2498 ? _T_10023 : _T_10030; // @[LoadQueue.scala 131:10:@13040.4]
  assign _T_10036 = 4'hd <= offsetQ_9; // @[LoadQueue.scala 131:81:@13043.4]
  assign _T_10037 = _T_6336 & _T_10036; // @[LoadQueue.scala 131:72:@13044.4]
  assign _T_10039 = offsetQ_9 < 4'hd; // @[LoadQueue.scala 132:33:@13045.4]
  assign _T_10042 = _T_10039 & _T_6345; // @[LoadQueue.scala 132:41:@13047.4]
  assign _T_10044 = _T_10042 == 1'h0; // @[LoadQueue.scala 132:9:@13048.4]
  assign storesToCheck_9_13 = _T_2498 ? _T_10037 : _T_10044; // @[LoadQueue.scala 131:10:@13049.4]
  assign _T_10050 = 4'he <= offsetQ_9; // @[LoadQueue.scala 131:81:@13052.4]
  assign _T_10051 = _T_6353 & _T_10050; // @[LoadQueue.scala 131:72:@13053.4]
  assign _T_10053 = offsetQ_9 < 4'he; // @[LoadQueue.scala 132:33:@13054.4]
  assign _T_10056 = _T_10053 & _T_6362; // @[LoadQueue.scala 132:41:@13056.4]
  assign _T_10058 = _T_10056 == 1'h0; // @[LoadQueue.scala 132:9:@13057.4]
  assign storesToCheck_9_14 = _T_2498 ? _T_10051 : _T_10058; // @[LoadQueue.scala 131:10:@13058.4]
  assign _T_10064 = 4'hf <= offsetQ_9; // @[LoadQueue.scala 131:81:@13061.4]
  assign storesToCheck_9_15 = _T_2498 ? _T_10064 : 1'h1; // @[LoadQueue.scala 131:10:@13067.4]
  assign storesToCheck_10_0 = _T_2528 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13109.4]
  assign _T_10114 = 4'h1 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13112.4]
  assign _T_10115 = _T_6132 & _T_10114; // @[LoadQueue.scala 131:72:@13113.4]
  assign _T_10117 = offsetQ_10 < 4'h1; // @[LoadQueue.scala 132:33:@13114.4]
  assign _T_10120 = _T_10117 & _T_6141; // @[LoadQueue.scala 132:41:@13116.4]
  assign _T_10122 = _T_10120 == 1'h0; // @[LoadQueue.scala 132:9:@13117.4]
  assign storesToCheck_10_1 = _T_2528 ? _T_10115 : _T_10122; // @[LoadQueue.scala 131:10:@13118.4]
  assign _T_10128 = 4'h2 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13121.4]
  assign _T_10129 = _T_6149 & _T_10128; // @[LoadQueue.scala 131:72:@13122.4]
  assign _T_10131 = offsetQ_10 < 4'h2; // @[LoadQueue.scala 132:33:@13123.4]
  assign _T_10134 = _T_10131 & _T_6158; // @[LoadQueue.scala 132:41:@13125.4]
  assign _T_10136 = _T_10134 == 1'h0; // @[LoadQueue.scala 132:9:@13126.4]
  assign storesToCheck_10_2 = _T_2528 ? _T_10129 : _T_10136; // @[LoadQueue.scala 131:10:@13127.4]
  assign _T_10142 = 4'h3 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13130.4]
  assign _T_10143 = _T_6166 & _T_10142; // @[LoadQueue.scala 131:72:@13131.4]
  assign _T_10145 = offsetQ_10 < 4'h3; // @[LoadQueue.scala 132:33:@13132.4]
  assign _T_10148 = _T_10145 & _T_6175; // @[LoadQueue.scala 132:41:@13134.4]
  assign _T_10150 = _T_10148 == 1'h0; // @[LoadQueue.scala 132:9:@13135.4]
  assign storesToCheck_10_3 = _T_2528 ? _T_10143 : _T_10150; // @[LoadQueue.scala 131:10:@13136.4]
  assign _T_10156 = 4'h4 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13139.4]
  assign _T_10157 = _T_6183 & _T_10156; // @[LoadQueue.scala 131:72:@13140.4]
  assign _T_10159 = offsetQ_10 < 4'h4; // @[LoadQueue.scala 132:33:@13141.4]
  assign _T_10162 = _T_10159 & _T_6192; // @[LoadQueue.scala 132:41:@13143.4]
  assign _T_10164 = _T_10162 == 1'h0; // @[LoadQueue.scala 132:9:@13144.4]
  assign storesToCheck_10_4 = _T_2528 ? _T_10157 : _T_10164; // @[LoadQueue.scala 131:10:@13145.4]
  assign _T_10170 = 4'h5 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13148.4]
  assign _T_10171 = _T_6200 & _T_10170; // @[LoadQueue.scala 131:72:@13149.4]
  assign _T_10173 = offsetQ_10 < 4'h5; // @[LoadQueue.scala 132:33:@13150.4]
  assign _T_10176 = _T_10173 & _T_6209; // @[LoadQueue.scala 132:41:@13152.4]
  assign _T_10178 = _T_10176 == 1'h0; // @[LoadQueue.scala 132:9:@13153.4]
  assign storesToCheck_10_5 = _T_2528 ? _T_10171 : _T_10178; // @[LoadQueue.scala 131:10:@13154.4]
  assign _T_10184 = 4'h6 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13157.4]
  assign _T_10185 = _T_6217 & _T_10184; // @[LoadQueue.scala 131:72:@13158.4]
  assign _T_10187 = offsetQ_10 < 4'h6; // @[LoadQueue.scala 132:33:@13159.4]
  assign _T_10190 = _T_10187 & _T_6226; // @[LoadQueue.scala 132:41:@13161.4]
  assign _T_10192 = _T_10190 == 1'h0; // @[LoadQueue.scala 132:9:@13162.4]
  assign storesToCheck_10_6 = _T_2528 ? _T_10185 : _T_10192; // @[LoadQueue.scala 131:10:@13163.4]
  assign _T_10198 = 4'h7 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13166.4]
  assign _T_10199 = _T_6234 & _T_10198; // @[LoadQueue.scala 131:72:@13167.4]
  assign _T_10201 = offsetQ_10 < 4'h7; // @[LoadQueue.scala 132:33:@13168.4]
  assign _T_10204 = _T_10201 & _T_6243; // @[LoadQueue.scala 132:41:@13170.4]
  assign _T_10206 = _T_10204 == 1'h0; // @[LoadQueue.scala 132:9:@13171.4]
  assign storesToCheck_10_7 = _T_2528 ? _T_10199 : _T_10206; // @[LoadQueue.scala 131:10:@13172.4]
  assign _T_10212 = 4'h8 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13175.4]
  assign _T_10213 = _T_6251 & _T_10212; // @[LoadQueue.scala 131:72:@13176.4]
  assign _T_10215 = offsetQ_10 < 4'h8; // @[LoadQueue.scala 132:33:@13177.4]
  assign _T_10218 = _T_10215 & _T_6260; // @[LoadQueue.scala 132:41:@13179.4]
  assign _T_10220 = _T_10218 == 1'h0; // @[LoadQueue.scala 132:9:@13180.4]
  assign storesToCheck_10_8 = _T_2528 ? _T_10213 : _T_10220; // @[LoadQueue.scala 131:10:@13181.4]
  assign _T_10226 = 4'h9 <= offsetQ_10; // @[LoadQueue.scala 131:81:@13184.4]
  assign _T_10227 = _T_6268 & _T_10226; // @[LoadQueue.scala 131:72:@13185.4]
  assign _T_10229 = offsetQ_10 < 4'h9; // @[LoadQueue.scala 132:33:@13186.4]
  assign _T_10232 = _T_10229 & _T_6277; // @[LoadQueue.scala 132:41:@13188.4]
  assign _T_10234 = _T_10232 == 1'h0; // @[LoadQueue.scala 132:9:@13189.4]
  assign storesToCheck_10_9 = _T_2528 ? _T_10227 : _T_10234; // @[LoadQueue.scala 131:10:@13190.4]
  assign _T_10240 = 4'ha <= offsetQ_10; // @[LoadQueue.scala 131:81:@13193.4]
  assign _T_10241 = _T_6285 & _T_10240; // @[LoadQueue.scala 131:72:@13194.4]
  assign _T_10243 = offsetQ_10 < 4'ha; // @[LoadQueue.scala 132:33:@13195.4]
  assign _T_10246 = _T_10243 & _T_6294; // @[LoadQueue.scala 132:41:@13197.4]
  assign _T_10248 = _T_10246 == 1'h0; // @[LoadQueue.scala 132:9:@13198.4]
  assign storesToCheck_10_10 = _T_2528 ? _T_10241 : _T_10248; // @[LoadQueue.scala 131:10:@13199.4]
  assign _T_10254 = 4'hb <= offsetQ_10; // @[LoadQueue.scala 131:81:@13202.4]
  assign _T_10255 = _T_6302 & _T_10254; // @[LoadQueue.scala 131:72:@13203.4]
  assign _T_10257 = offsetQ_10 < 4'hb; // @[LoadQueue.scala 132:33:@13204.4]
  assign _T_10260 = _T_10257 & _T_6311; // @[LoadQueue.scala 132:41:@13206.4]
  assign _T_10262 = _T_10260 == 1'h0; // @[LoadQueue.scala 132:9:@13207.4]
  assign storesToCheck_10_11 = _T_2528 ? _T_10255 : _T_10262; // @[LoadQueue.scala 131:10:@13208.4]
  assign _T_10268 = 4'hc <= offsetQ_10; // @[LoadQueue.scala 131:81:@13211.4]
  assign _T_10269 = _T_6319 & _T_10268; // @[LoadQueue.scala 131:72:@13212.4]
  assign _T_10271 = offsetQ_10 < 4'hc; // @[LoadQueue.scala 132:33:@13213.4]
  assign _T_10274 = _T_10271 & _T_6328; // @[LoadQueue.scala 132:41:@13215.4]
  assign _T_10276 = _T_10274 == 1'h0; // @[LoadQueue.scala 132:9:@13216.4]
  assign storesToCheck_10_12 = _T_2528 ? _T_10269 : _T_10276; // @[LoadQueue.scala 131:10:@13217.4]
  assign _T_10282 = 4'hd <= offsetQ_10; // @[LoadQueue.scala 131:81:@13220.4]
  assign _T_10283 = _T_6336 & _T_10282; // @[LoadQueue.scala 131:72:@13221.4]
  assign _T_10285 = offsetQ_10 < 4'hd; // @[LoadQueue.scala 132:33:@13222.4]
  assign _T_10288 = _T_10285 & _T_6345; // @[LoadQueue.scala 132:41:@13224.4]
  assign _T_10290 = _T_10288 == 1'h0; // @[LoadQueue.scala 132:9:@13225.4]
  assign storesToCheck_10_13 = _T_2528 ? _T_10283 : _T_10290; // @[LoadQueue.scala 131:10:@13226.4]
  assign _T_10296 = 4'he <= offsetQ_10; // @[LoadQueue.scala 131:81:@13229.4]
  assign _T_10297 = _T_6353 & _T_10296; // @[LoadQueue.scala 131:72:@13230.4]
  assign _T_10299 = offsetQ_10 < 4'he; // @[LoadQueue.scala 132:33:@13231.4]
  assign _T_10302 = _T_10299 & _T_6362; // @[LoadQueue.scala 132:41:@13233.4]
  assign _T_10304 = _T_10302 == 1'h0; // @[LoadQueue.scala 132:9:@13234.4]
  assign storesToCheck_10_14 = _T_2528 ? _T_10297 : _T_10304; // @[LoadQueue.scala 131:10:@13235.4]
  assign _T_10310 = 4'hf <= offsetQ_10; // @[LoadQueue.scala 131:81:@13238.4]
  assign storesToCheck_10_15 = _T_2528 ? _T_10310 : 1'h1; // @[LoadQueue.scala 131:10:@13244.4]
  assign storesToCheck_11_0 = _T_2558 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13286.4]
  assign _T_10360 = 4'h1 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13289.4]
  assign _T_10361 = _T_6132 & _T_10360; // @[LoadQueue.scala 131:72:@13290.4]
  assign _T_10363 = offsetQ_11 < 4'h1; // @[LoadQueue.scala 132:33:@13291.4]
  assign _T_10366 = _T_10363 & _T_6141; // @[LoadQueue.scala 132:41:@13293.4]
  assign _T_10368 = _T_10366 == 1'h0; // @[LoadQueue.scala 132:9:@13294.4]
  assign storesToCheck_11_1 = _T_2558 ? _T_10361 : _T_10368; // @[LoadQueue.scala 131:10:@13295.4]
  assign _T_10374 = 4'h2 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13298.4]
  assign _T_10375 = _T_6149 & _T_10374; // @[LoadQueue.scala 131:72:@13299.4]
  assign _T_10377 = offsetQ_11 < 4'h2; // @[LoadQueue.scala 132:33:@13300.4]
  assign _T_10380 = _T_10377 & _T_6158; // @[LoadQueue.scala 132:41:@13302.4]
  assign _T_10382 = _T_10380 == 1'h0; // @[LoadQueue.scala 132:9:@13303.4]
  assign storesToCheck_11_2 = _T_2558 ? _T_10375 : _T_10382; // @[LoadQueue.scala 131:10:@13304.4]
  assign _T_10388 = 4'h3 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13307.4]
  assign _T_10389 = _T_6166 & _T_10388; // @[LoadQueue.scala 131:72:@13308.4]
  assign _T_10391 = offsetQ_11 < 4'h3; // @[LoadQueue.scala 132:33:@13309.4]
  assign _T_10394 = _T_10391 & _T_6175; // @[LoadQueue.scala 132:41:@13311.4]
  assign _T_10396 = _T_10394 == 1'h0; // @[LoadQueue.scala 132:9:@13312.4]
  assign storesToCheck_11_3 = _T_2558 ? _T_10389 : _T_10396; // @[LoadQueue.scala 131:10:@13313.4]
  assign _T_10402 = 4'h4 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13316.4]
  assign _T_10403 = _T_6183 & _T_10402; // @[LoadQueue.scala 131:72:@13317.4]
  assign _T_10405 = offsetQ_11 < 4'h4; // @[LoadQueue.scala 132:33:@13318.4]
  assign _T_10408 = _T_10405 & _T_6192; // @[LoadQueue.scala 132:41:@13320.4]
  assign _T_10410 = _T_10408 == 1'h0; // @[LoadQueue.scala 132:9:@13321.4]
  assign storesToCheck_11_4 = _T_2558 ? _T_10403 : _T_10410; // @[LoadQueue.scala 131:10:@13322.4]
  assign _T_10416 = 4'h5 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13325.4]
  assign _T_10417 = _T_6200 & _T_10416; // @[LoadQueue.scala 131:72:@13326.4]
  assign _T_10419 = offsetQ_11 < 4'h5; // @[LoadQueue.scala 132:33:@13327.4]
  assign _T_10422 = _T_10419 & _T_6209; // @[LoadQueue.scala 132:41:@13329.4]
  assign _T_10424 = _T_10422 == 1'h0; // @[LoadQueue.scala 132:9:@13330.4]
  assign storesToCheck_11_5 = _T_2558 ? _T_10417 : _T_10424; // @[LoadQueue.scala 131:10:@13331.4]
  assign _T_10430 = 4'h6 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13334.4]
  assign _T_10431 = _T_6217 & _T_10430; // @[LoadQueue.scala 131:72:@13335.4]
  assign _T_10433 = offsetQ_11 < 4'h6; // @[LoadQueue.scala 132:33:@13336.4]
  assign _T_10436 = _T_10433 & _T_6226; // @[LoadQueue.scala 132:41:@13338.4]
  assign _T_10438 = _T_10436 == 1'h0; // @[LoadQueue.scala 132:9:@13339.4]
  assign storesToCheck_11_6 = _T_2558 ? _T_10431 : _T_10438; // @[LoadQueue.scala 131:10:@13340.4]
  assign _T_10444 = 4'h7 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13343.4]
  assign _T_10445 = _T_6234 & _T_10444; // @[LoadQueue.scala 131:72:@13344.4]
  assign _T_10447 = offsetQ_11 < 4'h7; // @[LoadQueue.scala 132:33:@13345.4]
  assign _T_10450 = _T_10447 & _T_6243; // @[LoadQueue.scala 132:41:@13347.4]
  assign _T_10452 = _T_10450 == 1'h0; // @[LoadQueue.scala 132:9:@13348.4]
  assign storesToCheck_11_7 = _T_2558 ? _T_10445 : _T_10452; // @[LoadQueue.scala 131:10:@13349.4]
  assign _T_10458 = 4'h8 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13352.4]
  assign _T_10459 = _T_6251 & _T_10458; // @[LoadQueue.scala 131:72:@13353.4]
  assign _T_10461 = offsetQ_11 < 4'h8; // @[LoadQueue.scala 132:33:@13354.4]
  assign _T_10464 = _T_10461 & _T_6260; // @[LoadQueue.scala 132:41:@13356.4]
  assign _T_10466 = _T_10464 == 1'h0; // @[LoadQueue.scala 132:9:@13357.4]
  assign storesToCheck_11_8 = _T_2558 ? _T_10459 : _T_10466; // @[LoadQueue.scala 131:10:@13358.4]
  assign _T_10472 = 4'h9 <= offsetQ_11; // @[LoadQueue.scala 131:81:@13361.4]
  assign _T_10473 = _T_6268 & _T_10472; // @[LoadQueue.scala 131:72:@13362.4]
  assign _T_10475 = offsetQ_11 < 4'h9; // @[LoadQueue.scala 132:33:@13363.4]
  assign _T_10478 = _T_10475 & _T_6277; // @[LoadQueue.scala 132:41:@13365.4]
  assign _T_10480 = _T_10478 == 1'h0; // @[LoadQueue.scala 132:9:@13366.4]
  assign storesToCheck_11_9 = _T_2558 ? _T_10473 : _T_10480; // @[LoadQueue.scala 131:10:@13367.4]
  assign _T_10486 = 4'ha <= offsetQ_11; // @[LoadQueue.scala 131:81:@13370.4]
  assign _T_10487 = _T_6285 & _T_10486; // @[LoadQueue.scala 131:72:@13371.4]
  assign _T_10489 = offsetQ_11 < 4'ha; // @[LoadQueue.scala 132:33:@13372.4]
  assign _T_10492 = _T_10489 & _T_6294; // @[LoadQueue.scala 132:41:@13374.4]
  assign _T_10494 = _T_10492 == 1'h0; // @[LoadQueue.scala 132:9:@13375.4]
  assign storesToCheck_11_10 = _T_2558 ? _T_10487 : _T_10494; // @[LoadQueue.scala 131:10:@13376.4]
  assign _T_10500 = 4'hb <= offsetQ_11; // @[LoadQueue.scala 131:81:@13379.4]
  assign _T_10501 = _T_6302 & _T_10500; // @[LoadQueue.scala 131:72:@13380.4]
  assign _T_10503 = offsetQ_11 < 4'hb; // @[LoadQueue.scala 132:33:@13381.4]
  assign _T_10506 = _T_10503 & _T_6311; // @[LoadQueue.scala 132:41:@13383.4]
  assign _T_10508 = _T_10506 == 1'h0; // @[LoadQueue.scala 132:9:@13384.4]
  assign storesToCheck_11_11 = _T_2558 ? _T_10501 : _T_10508; // @[LoadQueue.scala 131:10:@13385.4]
  assign _T_10514 = 4'hc <= offsetQ_11; // @[LoadQueue.scala 131:81:@13388.4]
  assign _T_10515 = _T_6319 & _T_10514; // @[LoadQueue.scala 131:72:@13389.4]
  assign _T_10517 = offsetQ_11 < 4'hc; // @[LoadQueue.scala 132:33:@13390.4]
  assign _T_10520 = _T_10517 & _T_6328; // @[LoadQueue.scala 132:41:@13392.4]
  assign _T_10522 = _T_10520 == 1'h0; // @[LoadQueue.scala 132:9:@13393.4]
  assign storesToCheck_11_12 = _T_2558 ? _T_10515 : _T_10522; // @[LoadQueue.scala 131:10:@13394.4]
  assign _T_10528 = 4'hd <= offsetQ_11; // @[LoadQueue.scala 131:81:@13397.4]
  assign _T_10529 = _T_6336 & _T_10528; // @[LoadQueue.scala 131:72:@13398.4]
  assign _T_10531 = offsetQ_11 < 4'hd; // @[LoadQueue.scala 132:33:@13399.4]
  assign _T_10534 = _T_10531 & _T_6345; // @[LoadQueue.scala 132:41:@13401.4]
  assign _T_10536 = _T_10534 == 1'h0; // @[LoadQueue.scala 132:9:@13402.4]
  assign storesToCheck_11_13 = _T_2558 ? _T_10529 : _T_10536; // @[LoadQueue.scala 131:10:@13403.4]
  assign _T_10542 = 4'he <= offsetQ_11; // @[LoadQueue.scala 131:81:@13406.4]
  assign _T_10543 = _T_6353 & _T_10542; // @[LoadQueue.scala 131:72:@13407.4]
  assign _T_10545 = offsetQ_11 < 4'he; // @[LoadQueue.scala 132:33:@13408.4]
  assign _T_10548 = _T_10545 & _T_6362; // @[LoadQueue.scala 132:41:@13410.4]
  assign _T_10550 = _T_10548 == 1'h0; // @[LoadQueue.scala 132:9:@13411.4]
  assign storesToCheck_11_14 = _T_2558 ? _T_10543 : _T_10550; // @[LoadQueue.scala 131:10:@13412.4]
  assign _T_10556 = 4'hf <= offsetQ_11; // @[LoadQueue.scala 131:81:@13415.4]
  assign storesToCheck_11_15 = _T_2558 ? _T_10556 : 1'h1; // @[LoadQueue.scala 131:10:@13421.4]
  assign storesToCheck_12_0 = _T_2588 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13463.4]
  assign _T_10606 = 4'h1 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13466.4]
  assign _T_10607 = _T_6132 & _T_10606; // @[LoadQueue.scala 131:72:@13467.4]
  assign _T_10609 = offsetQ_12 < 4'h1; // @[LoadQueue.scala 132:33:@13468.4]
  assign _T_10612 = _T_10609 & _T_6141; // @[LoadQueue.scala 132:41:@13470.4]
  assign _T_10614 = _T_10612 == 1'h0; // @[LoadQueue.scala 132:9:@13471.4]
  assign storesToCheck_12_1 = _T_2588 ? _T_10607 : _T_10614; // @[LoadQueue.scala 131:10:@13472.4]
  assign _T_10620 = 4'h2 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13475.4]
  assign _T_10621 = _T_6149 & _T_10620; // @[LoadQueue.scala 131:72:@13476.4]
  assign _T_10623 = offsetQ_12 < 4'h2; // @[LoadQueue.scala 132:33:@13477.4]
  assign _T_10626 = _T_10623 & _T_6158; // @[LoadQueue.scala 132:41:@13479.4]
  assign _T_10628 = _T_10626 == 1'h0; // @[LoadQueue.scala 132:9:@13480.4]
  assign storesToCheck_12_2 = _T_2588 ? _T_10621 : _T_10628; // @[LoadQueue.scala 131:10:@13481.4]
  assign _T_10634 = 4'h3 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13484.4]
  assign _T_10635 = _T_6166 & _T_10634; // @[LoadQueue.scala 131:72:@13485.4]
  assign _T_10637 = offsetQ_12 < 4'h3; // @[LoadQueue.scala 132:33:@13486.4]
  assign _T_10640 = _T_10637 & _T_6175; // @[LoadQueue.scala 132:41:@13488.4]
  assign _T_10642 = _T_10640 == 1'h0; // @[LoadQueue.scala 132:9:@13489.4]
  assign storesToCheck_12_3 = _T_2588 ? _T_10635 : _T_10642; // @[LoadQueue.scala 131:10:@13490.4]
  assign _T_10648 = 4'h4 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13493.4]
  assign _T_10649 = _T_6183 & _T_10648; // @[LoadQueue.scala 131:72:@13494.4]
  assign _T_10651 = offsetQ_12 < 4'h4; // @[LoadQueue.scala 132:33:@13495.4]
  assign _T_10654 = _T_10651 & _T_6192; // @[LoadQueue.scala 132:41:@13497.4]
  assign _T_10656 = _T_10654 == 1'h0; // @[LoadQueue.scala 132:9:@13498.4]
  assign storesToCheck_12_4 = _T_2588 ? _T_10649 : _T_10656; // @[LoadQueue.scala 131:10:@13499.4]
  assign _T_10662 = 4'h5 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13502.4]
  assign _T_10663 = _T_6200 & _T_10662; // @[LoadQueue.scala 131:72:@13503.4]
  assign _T_10665 = offsetQ_12 < 4'h5; // @[LoadQueue.scala 132:33:@13504.4]
  assign _T_10668 = _T_10665 & _T_6209; // @[LoadQueue.scala 132:41:@13506.4]
  assign _T_10670 = _T_10668 == 1'h0; // @[LoadQueue.scala 132:9:@13507.4]
  assign storesToCheck_12_5 = _T_2588 ? _T_10663 : _T_10670; // @[LoadQueue.scala 131:10:@13508.4]
  assign _T_10676 = 4'h6 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13511.4]
  assign _T_10677 = _T_6217 & _T_10676; // @[LoadQueue.scala 131:72:@13512.4]
  assign _T_10679 = offsetQ_12 < 4'h6; // @[LoadQueue.scala 132:33:@13513.4]
  assign _T_10682 = _T_10679 & _T_6226; // @[LoadQueue.scala 132:41:@13515.4]
  assign _T_10684 = _T_10682 == 1'h0; // @[LoadQueue.scala 132:9:@13516.4]
  assign storesToCheck_12_6 = _T_2588 ? _T_10677 : _T_10684; // @[LoadQueue.scala 131:10:@13517.4]
  assign _T_10690 = 4'h7 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13520.4]
  assign _T_10691 = _T_6234 & _T_10690; // @[LoadQueue.scala 131:72:@13521.4]
  assign _T_10693 = offsetQ_12 < 4'h7; // @[LoadQueue.scala 132:33:@13522.4]
  assign _T_10696 = _T_10693 & _T_6243; // @[LoadQueue.scala 132:41:@13524.4]
  assign _T_10698 = _T_10696 == 1'h0; // @[LoadQueue.scala 132:9:@13525.4]
  assign storesToCheck_12_7 = _T_2588 ? _T_10691 : _T_10698; // @[LoadQueue.scala 131:10:@13526.4]
  assign _T_10704 = 4'h8 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13529.4]
  assign _T_10705 = _T_6251 & _T_10704; // @[LoadQueue.scala 131:72:@13530.4]
  assign _T_10707 = offsetQ_12 < 4'h8; // @[LoadQueue.scala 132:33:@13531.4]
  assign _T_10710 = _T_10707 & _T_6260; // @[LoadQueue.scala 132:41:@13533.4]
  assign _T_10712 = _T_10710 == 1'h0; // @[LoadQueue.scala 132:9:@13534.4]
  assign storesToCheck_12_8 = _T_2588 ? _T_10705 : _T_10712; // @[LoadQueue.scala 131:10:@13535.4]
  assign _T_10718 = 4'h9 <= offsetQ_12; // @[LoadQueue.scala 131:81:@13538.4]
  assign _T_10719 = _T_6268 & _T_10718; // @[LoadQueue.scala 131:72:@13539.4]
  assign _T_10721 = offsetQ_12 < 4'h9; // @[LoadQueue.scala 132:33:@13540.4]
  assign _T_10724 = _T_10721 & _T_6277; // @[LoadQueue.scala 132:41:@13542.4]
  assign _T_10726 = _T_10724 == 1'h0; // @[LoadQueue.scala 132:9:@13543.4]
  assign storesToCheck_12_9 = _T_2588 ? _T_10719 : _T_10726; // @[LoadQueue.scala 131:10:@13544.4]
  assign _T_10732 = 4'ha <= offsetQ_12; // @[LoadQueue.scala 131:81:@13547.4]
  assign _T_10733 = _T_6285 & _T_10732; // @[LoadQueue.scala 131:72:@13548.4]
  assign _T_10735 = offsetQ_12 < 4'ha; // @[LoadQueue.scala 132:33:@13549.4]
  assign _T_10738 = _T_10735 & _T_6294; // @[LoadQueue.scala 132:41:@13551.4]
  assign _T_10740 = _T_10738 == 1'h0; // @[LoadQueue.scala 132:9:@13552.4]
  assign storesToCheck_12_10 = _T_2588 ? _T_10733 : _T_10740; // @[LoadQueue.scala 131:10:@13553.4]
  assign _T_10746 = 4'hb <= offsetQ_12; // @[LoadQueue.scala 131:81:@13556.4]
  assign _T_10747 = _T_6302 & _T_10746; // @[LoadQueue.scala 131:72:@13557.4]
  assign _T_10749 = offsetQ_12 < 4'hb; // @[LoadQueue.scala 132:33:@13558.4]
  assign _T_10752 = _T_10749 & _T_6311; // @[LoadQueue.scala 132:41:@13560.4]
  assign _T_10754 = _T_10752 == 1'h0; // @[LoadQueue.scala 132:9:@13561.4]
  assign storesToCheck_12_11 = _T_2588 ? _T_10747 : _T_10754; // @[LoadQueue.scala 131:10:@13562.4]
  assign _T_10760 = 4'hc <= offsetQ_12; // @[LoadQueue.scala 131:81:@13565.4]
  assign _T_10761 = _T_6319 & _T_10760; // @[LoadQueue.scala 131:72:@13566.4]
  assign _T_10763 = offsetQ_12 < 4'hc; // @[LoadQueue.scala 132:33:@13567.4]
  assign _T_10766 = _T_10763 & _T_6328; // @[LoadQueue.scala 132:41:@13569.4]
  assign _T_10768 = _T_10766 == 1'h0; // @[LoadQueue.scala 132:9:@13570.4]
  assign storesToCheck_12_12 = _T_2588 ? _T_10761 : _T_10768; // @[LoadQueue.scala 131:10:@13571.4]
  assign _T_10774 = 4'hd <= offsetQ_12; // @[LoadQueue.scala 131:81:@13574.4]
  assign _T_10775 = _T_6336 & _T_10774; // @[LoadQueue.scala 131:72:@13575.4]
  assign _T_10777 = offsetQ_12 < 4'hd; // @[LoadQueue.scala 132:33:@13576.4]
  assign _T_10780 = _T_10777 & _T_6345; // @[LoadQueue.scala 132:41:@13578.4]
  assign _T_10782 = _T_10780 == 1'h0; // @[LoadQueue.scala 132:9:@13579.4]
  assign storesToCheck_12_13 = _T_2588 ? _T_10775 : _T_10782; // @[LoadQueue.scala 131:10:@13580.4]
  assign _T_10788 = 4'he <= offsetQ_12; // @[LoadQueue.scala 131:81:@13583.4]
  assign _T_10789 = _T_6353 & _T_10788; // @[LoadQueue.scala 131:72:@13584.4]
  assign _T_10791 = offsetQ_12 < 4'he; // @[LoadQueue.scala 132:33:@13585.4]
  assign _T_10794 = _T_10791 & _T_6362; // @[LoadQueue.scala 132:41:@13587.4]
  assign _T_10796 = _T_10794 == 1'h0; // @[LoadQueue.scala 132:9:@13588.4]
  assign storesToCheck_12_14 = _T_2588 ? _T_10789 : _T_10796; // @[LoadQueue.scala 131:10:@13589.4]
  assign _T_10802 = 4'hf <= offsetQ_12; // @[LoadQueue.scala 131:81:@13592.4]
  assign storesToCheck_12_15 = _T_2588 ? _T_10802 : 1'h1; // @[LoadQueue.scala 131:10:@13598.4]
  assign storesToCheck_13_0 = _T_2618 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13640.4]
  assign _T_10852 = 4'h1 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13643.4]
  assign _T_10853 = _T_6132 & _T_10852; // @[LoadQueue.scala 131:72:@13644.4]
  assign _T_10855 = offsetQ_13 < 4'h1; // @[LoadQueue.scala 132:33:@13645.4]
  assign _T_10858 = _T_10855 & _T_6141; // @[LoadQueue.scala 132:41:@13647.4]
  assign _T_10860 = _T_10858 == 1'h0; // @[LoadQueue.scala 132:9:@13648.4]
  assign storesToCheck_13_1 = _T_2618 ? _T_10853 : _T_10860; // @[LoadQueue.scala 131:10:@13649.4]
  assign _T_10866 = 4'h2 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13652.4]
  assign _T_10867 = _T_6149 & _T_10866; // @[LoadQueue.scala 131:72:@13653.4]
  assign _T_10869 = offsetQ_13 < 4'h2; // @[LoadQueue.scala 132:33:@13654.4]
  assign _T_10872 = _T_10869 & _T_6158; // @[LoadQueue.scala 132:41:@13656.4]
  assign _T_10874 = _T_10872 == 1'h0; // @[LoadQueue.scala 132:9:@13657.4]
  assign storesToCheck_13_2 = _T_2618 ? _T_10867 : _T_10874; // @[LoadQueue.scala 131:10:@13658.4]
  assign _T_10880 = 4'h3 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13661.4]
  assign _T_10881 = _T_6166 & _T_10880; // @[LoadQueue.scala 131:72:@13662.4]
  assign _T_10883 = offsetQ_13 < 4'h3; // @[LoadQueue.scala 132:33:@13663.4]
  assign _T_10886 = _T_10883 & _T_6175; // @[LoadQueue.scala 132:41:@13665.4]
  assign _T_10888 = _T_10886 == 1'h0; // @[LoadQueue.scala 132:9:@13666.4]
  assign storesToCheck_13_3 = _T_2618 ? _T_10881 : _T_10888; // @[LoadQueue.scala 131:10:@13667.4]
  assign _T_10894 = 4'h4 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13670.4]
  assign _T_10895 = _T_6183 & _T_10894; // @[LoadQueue.scala 131:72:@13671.4]
  assign _T_10897 = offsetQ_13 < 4'h4; // @[LoadQueue.scala 132:33:@13672.4]
  assign _T_10900 = _T_10897 & _T_6192; // @[LoadQueue.scala 132:41:@13674.4]
  assign _T_10902 = _T_10900 == 1'h0; // @[LoadQueue.scala 132:9:@13675.4]
  assign storesToCheck_13_4 = _T_2618 ? _T_10895 : _T_10902; // @[LoadQueue.scala 131:10:@13676.4]
  assign _T_10908 = 4'h5 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13679.4]
  assign _T_10909 = _T_6200 & _T_10908; // @[LoadQueue.scala 131:72:@13680.4]
  assign _T_10911 = offsetQ_13 < 4'h5; // @[LoadQueue.scala 132:33:@13681.4]
  assign _T_10914 = _T_10911 & _T_6209; // @[LoadQueue.scala 132:41:@13683.4]
  assign _T_10916 = _T_10914 == 1'h0; // @[LoadQueue.scala 132:9:@13684.4]
  assign storesToCheck_13_5 = _T_2618 ? _T_10909 : _T_10916; // @[LoadQueue.scala 131:10:@13685.4]
  assign _T_10922 = 4'h6 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13688.4]
  assign _T_10923 = _T_6217 & _T_10922; // @[LoadQueue.scala 131:72:@13689.4]
  assign _T_10925 = offsetQ_13 < 4'h6; // @[LoadQueue.scala 132:33:@13690.4]
  assign _T_10928 = _T_10925 & _T_6226; // @[LoadQueue.scala 132:41:@13692.4]
  assign _T_10930 = _T_10928 == 1'h0; // @[LoadQueue.scala 132:9:@13693.4]
  assign storesToCheck_13_6 = _T_2618 ? _T_10923 : _T_10930; // @[LoadQueue.scala 131:10:@13694.4]
  assign _T_10936 = 4'h7 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13697.4]
  assign _T_10937 = _T_6234 & _T_10936; // @[LoadQueue.scala 131:72:@13698.4]
  assign _T_10939 = offsetQ_13 < 4'h7; // @[LoadQueue.scala 132:33:@13699.4]
  assign _T_10942 = _T_10939 & _T_6243; // @[LoadQueue.scala 132:41:@13701.4]
  assign _T_10944 = _T_10942 == 1'h0; // @[LoadQueue.scala 132:9:@13702.4]
  assign storesToCheck_13_7 = _T_2618 ? _T_10937 : _T_10944; // @[LoadQueue.scala 131:10:@13703.4]
  assign _T_10950 = 4'h8 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13706.4]
  assign _T_10951 = _T_6251 & _T_10950; // @[LoadQueue.scala 131:72:@13707.4]
  assign _T_10953 = offsetQ_13 < 4'h8; // @[LoadQueue.scala 132:33:@13708.4]
  assign _T_10956 = _T_10953 & _T_6260; // @[LoadQueue.scala 132:41:@13710.4]
  assign _T_10958 = _T_10956 == 1'h0; // @[LoadQueue.scala 132:9:@13711.4]
  assign storesToCheck_13_8 = _T_2618 ? _T_10951 : _T_10958; // @[LoadQueue.scala 131:10:@13712.4]
  assign _T_10964 = 4'h9 <= offsetQ_13; // @[LoadQueue.scala 131:81:@13715.4]
  assign _T_10965 = _T_6268 & _T_10964; // @[LoadQueue.scala 131:72:@13716.4]
  assign _T_10967 = offsetQ_13 < 4'h9; // @[LoadQueue.scala 132:33:@13717.4]
  assign _T_10970 = _T_10967 & _T_6277; // @[LoadQueue.scala 132:41:@13719.4]
  assign _T_10972 = _T_10970 == 1'h0; // @[LoadQueue.scala 132:9:@13720.4]
  assign storesToCheck_13_9 = _T_2618 ? _T_10965 : _T_10972; // @[LoadQueue.scala 131:10:@13721.4]
  assign _T_10978 = 4'ha <= offsetQ_13; // @[LoadQueue.scala 131:81:@13724.4]
  assign _T_10979 = _T_6285 & _T_10978; // @[LoadQueue.scala 131:72:@13725.4]
  assign _T_10981 = offsetQ_13 < 4'ha; // @[LoadQueue.scala 132:33:@13726.4]
  assign _T_10984 = _T_10981 & _T_6294; // @[LoadQueue.scala 132:41:@13728.4]
  assign _T_10986 = _T_10984 == 1'h0; // @[LoadQueue.scala 132:9:@13729.4]
  assign storesToCheck_13_10 = _T_2618 ? _T_10979 : _T_10986; // @[LoadQueue.scala 131:10:@13730.4]
  assign _T_10992 = 4'hb <= offsetQ_13; // @[LoadQueue.scala 131:81:@13733.4]
  assign _T_10993 = _T_6302 & _T_10992; // @[LoadQueue.scala 131:72:@13734.4]
  assign _T_10995 = offsetQ_13 < 4'hb; // @[LoadQueue.scala 132:33:@13735.4]
  assign _T_10998 = _T_10995 & _T_6311; // @[LoadQueue.scala 132:41:@13737.4]
  assign _T_11000 = _T_10998 == 1'h0; // @[LoadQueue.scala 132:9:@13738.4]
  assign storesToCheck_13_11 = _T_2618 ? _T_10993 : _T_11000; // @[LoadQueue.scala 131:10:@13739.4]
  assign _T_11006 = 4'hc <= offsetQ_13; // @[LoadQueue.scala 131:81:@13742.4]
  assign _T_11007 = _T_6319 & _T_11006; // @[LoadQueue.scala 131:72:@13743.4]
  assign _T_11009 = offsetQ_13 < 4'hc; // @[LoadQueue.scala 132:33:@13744.4]
  assign _T_11012 = _T_11009 & _T_6328; // @[LoadQueue.scala 132:41:@13746.4]
  assign _T_11014 = _T_11012 == 1'h0; // @[LoadQueue.scala 132:9:@13747.4]
  assign storesToCheck_13_12 = _T_2618 ? _T_11007 : _T_11014; // @[LoadQueue.scala 131:10:@13748.4]
  assign _T_11020 = 4'hd <= offsetQ_13; // @[LoadQueue.scala 131:81:@13751.4]
  assign _T_11021 = _T_6336 & _T_11020; // @[LoadQueue.scala 131:72:@13752.4]
  assign _T_11023 = offsetQ_13 < 4'hd; // @[LoadQueue.scala 132:33:@13753.4]
  assign _T_11026 = _T_11023 & _T_6345; // @[LoadQueue.scala 132:41:@13755.4]
  assign _T_11028 = _T_11026 == 1'h0; // @[LoadQueue.scala 132:9:@13756.4]
  assign storesToCheck_13_13 = _T_2618 ? _T_11021 : _T_11028; // @[LoadQueue.scala 131:10:@13757.4]
  assign _T_11034 = 4'he <= offsetQ_13; // @[LoadQueue.scala 131:81:@13760.4]
  assign _T_11035 = _T_6353 & _T_11034; // @[LoadQueue.scala 131:72:@13761.4]
  assign _T_11037 = offsetQ_13 < 4'he; // @[LoadQueue.scala 132:33:@13762.4]
  assign _T_11040 = _T_11037 & _T_6362; // @[LoadQueue.scala 132:41:@13764.4]
  assign _T_11042 = _T_11040 == 1'h0; // @[LoadQueue.scala 132:9:@13765.4]
  assign storesToCheck_13_14 = _T_2618 ? _T_11035 : _T_11042; // @[LoadQueue.scala 131:10:@13766.4]
  assign _T_11048 = 4'hf <= offsetQ_13; // @[LoadQueue.scala 131:81:@13769.4]
  assign storesToCheck_13_15 = _T_2618 ? _T_11048 : 1'h1; // @[LoadQueue.scala 131:10:@13775.4]
  assign storesToCheck_14_0 = _T_2648 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13817.4]
  assign _T_11098 = 4'h1 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13820.4]
  assign _T_11099 = _T_6132 & _T_11098; // @[LoadQueue.scala 131:72:@13821.4]
  assign _T_11101 = offsetQ_14 < 4'h1; // @[LoadQueue.scala 132:33:@13822.4]
  assign _T_11104 = _T_11101 & _T_6141; // @[LoadQueue.scala 132:41:@13824.4]
  assign _T_11106 = _T_11104 == 1'h0; // @[LoadQueue.scala 132:9:@13825.4]
  assign storesToCheck_14_1 = _T_2648 ? _T_11099 : _T_11106; // @[LoadQueue.scala 131:10:@13826.4]
  assign _T_11112 = 4'h2 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13829.4]
  assign _T_11113 = _T_6149 & _T_11112; // @[LoadQueue.scala 131:72:@13830.4]
  assign _T_11115 = offsetQ_14 < 4'h2; // @[LoadQueue.scala 132:33:@13831.4]
  assign _T_11118 = _T_11115 & _T_6158; // @[LoadQueue.scala 132:41:@13833.4]
  assign _T_11120 = _T_11118 == 1'h0; // @[LoadQueue.scala 132:9:@13834.4]
  assign storesToCheck_14_2 = _T_2648 ? _T_11113 : _T_11120; // @[LoadQueue.scala 131:10:@13835.4]
  assign _T_11126 = 4'h3 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13838.4]
  assign _T_11127 = _T_6166 & _T_11126; // @[LoadQueue.scala 131:72:@13839.4]
  assign _T_11129 = offsetQ_14 < 4'h3; // @[LoadQueue.scala 132:33:@13840.4]
  assign _T_11132 = _T_11129 & _T_6175; // @[LoadQueue.scala 132:41:@13842.4]
  assign _T_11134 = _T_11132 == 1'h0; // @[LoadQueue.scala 132:9:@13843.4]
  assign storesToCheck_14_3 = _T_2648 ? _T_11127 : _T_11134; // @[LoadQueue.scala 131:10:@13844.4]
  assign _T_11140 = 4'h4 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13847.4]
  assign _T_11141 = _T_6183 & _T_11140; // @[LoadQueue.scala 131:72:@13848.4]
  assign _T_11143 = offsetQ_14 < 4'h4; // @[LoadQueue.scala 132:33:@13849.4]
  assign _T_11146 = _T_11143 & _T_6192; // @[LoadQueue.scala 132:41:@13851.4]
  assign _T_11148 = _T_11146 == 1'h0; // @[LoadQueue.scala 132:9:@13852.4]
  assign storesToCheck_14_4 = _T_2648 ? _T_11141 : _T_11148; // @[LoadQueue.scala 131:10:@13853.4]
  assign _T_11154 = 4'h5 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13856.4]
  assign _T_11155 = _T_6200 & _T_11154; // @[LoadQueue.scala 131:72:@13857.4]
  assign _T_11157 = offsetQ_14 < 4'h5; // @[LoadQueue.scala 132:33:@13858.4]
  assign _T_11160 = _T_11157 & _T_6209; // @[LoadQueue.scala 132:41:@13860.4]
  assign _T_11162 = _T_11160 == 1'h0; // @[LoadQueue.scala 132:9:@13861.4]
  assign storesToCheck_14_5 = _T_2648 ? _T_11155 : _T_11162; // @[LoadQueue.scala 131:10:@13862.4]
  assign _T_11168 = 4'h6 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13865.4]
  assign _T_11169 = _T_6217 & _T_11168; // @[LoadQueue.scala 131:72:@13866.4]
  assign _T_11171 = offsetQ_14 < 4'h6; // @[LoadQueue.scala 132:33:@13867.4]
  assign _T_11174 = _T_11171 & _T_6226; // @[LoadQueue.scala 132:41:@13869.4]
  assign _T_11176 = _T_11174 == 1'h0; // @[LoadQueue.scala 132:9:@13870.4]
  assign storesToCheck_14_6 = _T_2648 ? _T_11169 : _T_11176; // @[LoadQueue.scala 131:10:@13871.4]
  assign _T_11182 = 4'h7 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13874.4]
  assign _T_11183 = _T_6234 & _T_11182; // @[LoadQueue.scala 131:72:@13875.4]
  assign _T_11185 = offsetQ_14 < 4'h7; // @[LoadQueue.scala 132:33:@13876.4]
  assign _T_11188 = _T_11185 & _T_6243; // @[LoadQueue.scala 132:41:@13878.4]
  assign _T_11190 = _T_11188 == 1'h0; // @[LoadQueue.scala 132:9:@13879.4]
  assign storesToCheck_14_7 = _T_2648 ? _T_11183 : _T_11190; // @[LoadQueue.scala 131:10:@13880.4]
  assign _T_11196 = 4'h8 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13883.4]
  assign _T_11197 = _T_6251 & _T_11196; // @[LoadQueue.scala 131:72:@13884.4]
  assign _T_11199 = offsetQ_14 < 4'h8; // @[LoadQueue.scala 132:33:@13885.4]
  assign _T_11202 = _T_11199 & _T_6260; // @[LoadQueue.scala 132:41:@13887.4]
  assign _T_11204 = _T_11202 == 1'h0; // @[LoadQueue.scala 132:9:@13888.4]
  assign storesToCheck_14_8 = _T_2648 ? _T_11197 : _T_11204; // @[LoadQueue.scala 131:10:@13889.4]
  assign _T_11210 = 4'h9 <= offsetQ_14; // @[LoadQueue.scala 131:81:@13892.4]
  assign _T_11211 = _T_6268 & _T_11210; // @[LoadQueue.scala 131:72:@13893.4]
  assign _T_11213 = offsetQ_14 < 4'h9; // @[LoadQueue.scala 132:33:@13894.4]
  assign _T_11216 = _T_11213 & _T_6277; // @[LoadQueue.scala 132:41:@13896.4]
  assign _T_11218 = _T_11216 == 1'h0; // @[LoadQueue.scala 132:9:@13897.4]
  assign storesToCheck_14_9 = _T_2648 ? _T_11211 : _T_11218; // @[LoadQueue.scala 131:10:@13898.4]
  assign _T_11224 = 4'ha <= offsetQ_14; // @[LoadQueue.scala 131:81:@13901.4]
  assign _T_11225 = _T_6285 & _T_11224; // @[LoadQueue.scala 131:72:@13902.4]
  assign _T_11227 = offsetQ_14 < 4'ha; // @[LoadQueue.scala 132:33:@13903.4]
  assign _T_11230 = _T_11227 & _T_6294; // @[LoadQueue.scala 132:41:@13905.4]
  assign _T_11232 = _T_11230 == 1'h0; // @[LoadQueue.scala 132:9:@13906.4]
  assign storesToCheck_14_10 = _T_2648 ? _T_11225 : _T_11232; // @[LoadQueue.scala 131:10:@13907.4]
  assign _T_11238 = 4'hb <= offsetQ_14; // @[LoadQueue.scala 131:81:@13910.4]
  assign _T_11239 = _T_6302 & _T_11238; // @[LoadQueue.scala 131:72:@13911.4]
  assign _T_11241 = offsetQ_14 < 4'hb; // @[LoadQueue.scala 132:33:@13912.4]
  assign _T_11244 = _T_11241 & _T_6311; // @[LoadQueue.scala 132:41:@13914.4]
  assign _T_11246 = _T_11244 == 1'h0; // @[LoadQueue.scala 132:9:@13915.4]
  assign storesToCheck_14_11 = _T_2648 ? _T_11239 : _T_11246; // @[LoadQueue.scala 131:10:@13916.4]
  assign _T_11252 = 4'hc <= offsetQ_14; // @[LoadQueue.scala 131:81:@13919.4]
  assign _T_11253 = _T_6319 & _T_11252; // @[LoadQueue.scala 131:72:@13920.4]
  assign _T_11255 = offsetQ_14 < 4'hc; // @[LoadQueue.scala 132:33:@13921.4]
  assign _T_11258 = _T_11255 & _T_6328; // @[LoadQueue.scala 132:41:@13923.4]
  assign _T_11260 = _T_11258 == 1'h0; // @[LoadQueue.scala 132:9:@13924.4]
  assign storesToCheck_14_12 = _T_2648 ? _T_11253 : _T_11260; // @[LoadQueue.scala 131:10:@13925.4]
  assign _T_11266 = 4'hd <= offsetQ_14; // @[LoadQueue.scala 131:81:@13928.4]
  assign _T_11267 = _T_6336 & _T_11266; // @[LoadQueue.scala 131:72:@13929.4]
  assign _T_11269 = offsetQ_14 < 4'hd; // @[LoadQueue.scala 132:33:@13930.4]
  assign _T_11272 = _T_11269 & _T_6345; // @[LoadQueue.scala 132:41:@13932.4]
  assign _T_11274 = _T_11272 == 1'h0; // @[LoadQueue.scala 132:9:@13933.4]
  assign storesToCheck_14_13 = _T_2648 ? _T_11267 : _T_11274; // @[LoadQueue.scala 131:10:@13934.4]
  assign _T_11280 = 4'he <= offsetQ_14; // @[LoadQueue.scala 131:81:@13937.4]
  assign _T_11281 = _T_6353 & _T_11280; // @[LoadQueue.scala 131:72:@13938.4]
  assign _T_11283 = offsetQ_14 < 4'he; // @[LoadQueue.scala 132:33:@13939.4]
  assign _T_11286 = _T_11283 & _T_6362; // @[LoadQueue.scala 132:41:@13941.4]
  assign _T_11288 = _T_11286 == 1'h0; // @[LoadQueue.scala 132:9:@13942.4]
  assign storesToCheck_14_14 = _T_2648 ? _T_11281 : _T_11288; // @[LoadQueue.scala 131:10:@13943.4]
  assign _T_11294 = 4'hf <= offsetQ_14; // @[LoadQueue.scala 131:81:@13946.4]
  assign storesToCheck_14_15 = _T_2648 ? _T_11294 : 1'h1; // @[LoadQueue.scala 131:10:@13952.4]
  assign storesToCheck_15_0 = _T_2678 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@13994.4]
  assign _T_11344 = 4'h1 <= offsetQ_15; // @[LoadQueue.scala 131:81:@13997.4]
  assign _T_11345 = _T_6132 & _T_11344; // @[LoadQueue.scala 131:72:@13998.4]
  assign _T_11347 = offsetQ_15 < 4'h1; // @[LoadQueue.scala 132:33:@13999.4]
  assign _T_11350 = _T_11347 & _T_6141; // @[LoadQueue.scala 132:41:@14001.4]
  assign _T_11352 = _T_11350 == 1'h0; // @[LoadQueue.scala 132:9:@14002.4]
  assign storesToCheck_15_1 = _T_2678 ? _T_11345 : _T_11352; // @[LoadQueue.scala 131:10:@14003.4]
  assign _T_11358 = 4'h2 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14006.4]
  assign _T_11359 = _T_6149 & _T_11358; // @[LoadQueue.scala 131:72:@14007.4]
  assign _T_11361 = offsetQ_15 < 4'h2; // @[LoadQueue.scala 132:33:@14008.4]
  assign _T_11364 = _T_11361 & _T_6158; // @[LoadQueue.scala 132:41:@14010.4]
  assign _T_11366 = _T_11364 == 1'h0; // @[LoadQueue.scala 132:9:@14011.4]
  assign storesToCheck_15_2 = _T_2678 ? _T_11359 : _T_11366; // @[LoadQueue.scala 131:10:@14012.4]
  assign _T_11372 = 4'h3 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14015.4]
  assign _T_11373 = _T_6166 & _T_11372; // @[LoadQueue.scala 131:72:@14016.4]
  assign _T_11375 = offsetQ_15 < 4'h3; // @[LoadQueue.scala 132:33:@14017.4]
  assign _T_11378 = _T_11375 & _T_6175; // @[LoadQueue.scala 132:41:@14019.4]
  assign _T_11380 = _T_11378 == 1'h0; // @[LoadQueue.scala 132:9:@14020.4]
  assign storesToCheck_15_3 = _T_2678 ? _T_11373 : _T_11380; // @[LoadQueue.scala 131:10:@14021.4]
  assign _T_11386 = 4'h4 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14024.4]
  assign _T_11387 = _T_6183 & _T_11386; // @[LoadQueue.scala 131:72:@14025.4]
  assign _T_11389 = offsetQ_15 < 4'h4; // @[LoadQueue.scala 132:33:@14026.4]
  assign _T_11392 = _T_11389 & _T_6192; // @[LoadQueue.scala 132:41:@14028.4]
  assign _T_11394 = _T_11392 == 1'h0; // @[LoadQueue.scala 132:9:@14029.4]
  assign storesToCheck_15_4 = _T_2678 ? _T_11387 : _T_11394; // @[LoadQueue.scala 131:10:@14030.4]
  assign _T_11400 = 4'h5 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14033.4]
  assign _T_11401 = _T_6200 & _T_11400; // @[LoadQueue.scala 131:72:@14034.4]
  assign _T_11403 = offsetQ_15 < 4'h5; // @[LoadQueue.scala 132:33:@14035.4]
  assign _T_11406 = _T_11403 & _T_6209; // @[LoadQueue.scala 132:41:@14037.4]
  assign _T_11408 = _T_11406 == 1'h0; // @[LoadQueue.scala 132:9:@14038.4]
  assign storesToCheck_15_5 = _T_2678 ? _T_11401 : _T_11408; // @[LoadQueue.scala 131:10:@14039.4]
  assign _T_11414 = 4'h6 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14042.4]
  assign _T_11415 = _T_6217 & _T_11414; // @[LoadQueue.scala 131:72:@14043.4]
  assign _T_11417 = offsetQ_15 < 4'h6; // @[LoadQueue.scala 132:33:@14044.4]
  assign _T_11420 = _T_11417 & _T_6226; // @[LoadQueue.scala 132:41:@14046.4]
  assign _T_11422 = _T_11420 == 1'h0; // @[LoadQueue.scala 132:9:@14047.4]
  assign storesToCheck_15_6 = _T_2678 ? _T_11415 : _T_11422; // @[LoadQueue.scala 131:10:@14048.4]
  assign _T_11428 = 4'h7 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14051.4]
  assign _T_11429 = _T_6234 & _T_11428; // @[LoadQueue.scala 131:72:@14052.4]
  assign _T_11431 = offsetQ_15 < 4'h7; // @[LoadQueue.scala 132:33:@14053.4]
  assign _T_11434 = _T_11431 & _T_6243; // @[LoadQueue.scala 132:41:@14055.4]
  assign _T_11436 = _T_11434 == 1'h0; // @[LoadQueue.scala 132:9:@14056.4]
  assign storesToCheck_15_7 = _T_2678 ? _T_11429 : _T_11436; // @[LoadQueue.scala 131:10:@14057.4]
  assign _T_11442 = 4'h8 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14060.4]
  assign _T_11443 = _T_6251 & _T_11442; // @[LoadQueue.scala 131:72:@14061.4]
  assign _T_11445 = offsetQ_15 < 4'h8; // @[LoadQueue.scala 132:33:@14062.4]
  assign _T_11448 = _T_11445 & _T_6260; // @[LoadQueue.scala 132:41:@14064.4]
  assign _T_11450 = _T_11448 == 1'h0; // @[LoadQueue.scala 132:9:@14065.4]
  assign storesToCheck_15_8 = _T_2678 ? _T_11443 : _T_11450; // @[LoadQueue.scala 131:10:@14066.4]
  assign _T_11456 = 4'h9 <= offsetQ_15; // @[LoadQueue.scala 131:81:@14069.4]
  assign _T_11457 = _T_6268 & _T_11456; // @[LoadQueue.scala 131:72:@14070.4]
  assign _T_11459 = offsetQ_15 < 4'h9; // @[LoadQueue.scala 132:33:@14071.4]
  assign _T_11462 = _T_11459 & _T_6277; // @[LoadQueue.scala 132:41:@14073.4]
  assign _T_11464 = _T_11462 == 1'h0; // @[LoadQueue.scala 132:9:@14074.4]
  assign storesToCheck_15_9 = _T_2678 ? _T_11457 : _T_11464; // @[LoadQueue.scala 131:10:@14075.4]
  assign _T_11470 = 4'ha <= offsetQ_15; // @[LoadQueue.scala 131:81:@14078.4]
  assign _T_11471 = _T_6285 & _T_11470; // @[LoadQueue.scala 131:72:@14079.4]
  assign _T_11473 = offsetQ_15 < 4'ha; // @[LoadQueue.scala 132:33:@14080.4]
  assign _T_11476 = _T_11473 & _T_6294; // @[LoadQueue.scala 132:41:@14082.4]
  assign _T_11478 = _T_11476 == 1'h0; // @[LoadQueue.scala 132:9:@14083.4]
  assign storesToCheck_15_10 = _T_2678 ? _T_11471 : _T_11478; // @[LoadQueue.scala 131:10:@14084.4]
  assign _T_11484 = 4'hb <= offsetQ_15; // @[LoadQueue.scala 131:81:@14087.4]
  assign _T_11485 = _T_6302 & _T_11484; // @[LoadQueue.scala 131:72:@14088.4]
  assign _T_11487 = offsetQ_15 < 4'hb; // @[LoadQueue.scala 132:33:@14089.4]
  assign _T_11490 = _T_11487 & _T_6311; // @[LoadQueue.scala 132:41:@14091.4]
  assign _T_11492 = _T_11490 == 1'h0; // @[LoadQueue.scala 132:9:@14092.4]
  assign storesToCheck_15_11 = _T_2678 ? _T_11485 : _T_11492; // @[LoadQueue.scala 131:10:@14093.4]
  assign _T_11498 = 4'hc <= offsetQ_15; // @[LoadQueue.scala 131:81:@14096.4]
  assign _T_11499 = _T_6319 & _T_11498; // @[LoadQueue.scala 131:72:@14097.4]
  assign _T_11501 = offsetQ_15 < 4'hc; // @[LoadQueue.scala 132:33:@14098.4]
  assign _T_11504 = _T_11501 & _T_6328; // @[LoadQueue.scala 132:41:@14100.4]
  assign _T_11506 = _T_11504 == 1'h0; // @[LoadQueue.scala 132:9:@14101.4]
  assign storesToCheck_15_12 = _T_2678 ? _T_11499 : _T_11506; // @[LoadQueue.scala 131:10:@14102.4]
  assign _T_11512 = 4'hd <= offsetQ_15; // @[LoadQueue.scala 131:81:@14105.4]
  assign _T_11513 = _T_6336 & _T_11512; // @[LoadQueue.scala 131:72:@14106.4]
  assign _T_11515 = offsetQ_15 < 4'hd; // @[LoadQueue.scala 132:33:@14107.4]
  assign _T_11518 = _T_11515 & _T_6345; // @[LoadQueue.scala 132:41:@14109.4]
  assign _T_11520 = _T_11518 == 1'h0; // @[LoadQueue.scala 132:9:@14110.4]
  assign storesToCheck_15_13 = _T_2678 ? _T_11513 : _T_11520; // @[LoadQueue.scala 131:10:@14111.4]
  assign _T_11526 = 4'he <= offsetQ_15; // @[LoadQueue.scala 131:81:@14114.4]
  assign _T_11527 = _T_6353 & _T_11526; // @[LoadQueue.scala 131:72:@14115.4]
  assign _T_11529 = offsetQ_15 < 4'he; // @[LoadQueue.scala 132:33:@14116.4]
  assign _T_11532 = _T_11529 & _T_6362; // @[LoadQueue.scala 132:41:@14118.4]
  assign _T_11534 = _T_11532 == 1'h0; // @[LoadQueue.scala 132:9:@14119.4]
  assign storesToCheck_15_14 = _T_2678 ? _T_11527 : _T_11534; // @[LoadQueue.scala 131:10:@14120.4]
  assign _T_11540 = 4'hf <= offsetQ_15; // @[LoadQueue.scala 131:81:@14123.4]
  assign storesToCheck_15_15 = _T_2678 ? _T_11540 : 1'h1; // @[LoadQueue.scala 131:10:@14129.4]
  assign _T_12802 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14164.4]
  assign entriesToCheck_0_0 = _T_12802 & checkBits_0; // @[LoadQueue.scala 141:26:@14165.4]
  assign _T_12804 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14166.4]
  assign entriesToCheck_0_1 = _T_12804 & checkBits_0; // @[LoadQueue.scala 141:26:@14167.4]
  assign _T_12806 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14168.4]
  assign entriesToCheck_0_2 = _T_12806 & checkBits_0; // @[LoadQueue.scala 141:26:@14169.4]
  assign _T_12808 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14170.4]
  assign entriesToCheck_0_3 = _T_12808 & checkBits_0; // @[LoadQueue.scala 141:26:@14171.4]
  assign _T_12810 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14172.4]
  assign entriesToCheck_0_4 = _T_12810 & checkBits_0; // @[LoadQueue.scala 141:26:@14173.4]
  assign _T_12812 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14174.4]
  assign entriesToCheck_0_5 = _T_12812 & checkBits_0; // @[LoadQueue.scala 141:26:@14175.4]
  assign _T_12814 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14176.4]
  assign entriesToCheck_0_6 = _T_12814 & checkBits_0; // @[LoadQueue.scala 141:26:@14177.4]
  assign _T_12816 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14178.4]
  assign entriesToCheck_0_7 = _T_12816 & checkBits_0; // @[LoadQueue.scala 141:26:@14179.4]
  assign _T_12818 = storesToCheck_0_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14180.4]
  assign entriesToCheck_0_8 = _T_12818 & checkBits_0; // @[LoadQueue.scala 141:26:@14181.4]
  assign _T_12820 = storesToCheck_0_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14182.4]
  assign entriesToCheck_0_9 = _T_12820 & checkBits_0; // @[LoadQueue.scala 141:26:@14183.4]
  assign _T_12822 = storesToCheck_0_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14184.4]
  assign entriesToCheck_0_10 = _T_12822 & checkBits_0; // @[LoadQueue.scala 141:26:@14185.4]
  assign _T_12824 = storesToCheck_0_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14186.4]
  assign entriesToCheck_0_11 = _T_12824 & checkBits_0; // @[LoadQueue.scala 141:26:@14187.4]
  assign _T_12826 = storesToCheck_0_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14188.4]
  assign entriesToCheck_0_12 = _T_12826 & checkBits_0; // @[LoadQueue.scala 141:26:@14189.4]
  assign _T_12828 = storesToCheck_0_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14190.4]
  assign entriesToCheck_0_13 = _T_12828 & checkBits_0; // @[LoadQueue.scala 141:26:@14191.4]
  assign _T_12830 = storesToCheck_0_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14192.4]
  assign entriesToCheck_0_14 = _T_12830 & checkBits_0; // @[LoadQueue.scala 141:26:@14193.4]
  assign _T_12832 = storesToCheck_0_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14194.4]
  assign entriesToCheck_0_15 = _T_12832 & checkBits_0; // @[LoadQueue.scala 141:26:@14195.4]
  assign _T_12834 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14212.4]
  assign entriesToCheck_1_0 = _T_12834 & checkBits_1; // @[LoadQueue.scala 141:26:@14213.4]
  assign _T_12836 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14214.4]
  assign entriesToCheck_1_1 = _T_12836 & checkBits_1; // @[LoadQueue.scala 141:26:@14215.4]
  assign _T_12838 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14216.4]
  assign entriesToCheck_1_2 = _T_12838 & checkBits_1; // @[LoadQueue.scala 141:26:@14217.4]
  assign _T_12840 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14218.4]
  assign entriesToCheck_1_3 = _T_12840 & checkBits_1; // @[LoadQueue.scala 141:26:@14219.4]
  assign _T_12842 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14220.4]
  assign entriesToCheck_1_4 = _T_12842 & checkBits_1; // @[LoadQueue.scala 141:26:@14221.4]
  assign _T_12844 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14222.4]
  assign entriesToCheck_1_5 = _T_12844 & checkBits_1; // @[LoadQueue.scala 141:26:@14223.4]
  assign _T_12846 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14224.4]
  assign entriesToCheck_1_6 = _T_12846 & checkBits_1; // @[LoadQueue.scala 141:26:@14225.4]
  assign _T_12848 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14226.4]
  assign entriesToCheck_1_7 = _T_12848 & checkBits_1; // @[LoadQueue.scala 141:26:@14227.4]
  assign _T_12850 = storesToCheck_1_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14228.4]
  assign entriesToCheck_1_8 = _T_12850 & checkBits_1; // @[LoadQueue.scala 141:26:@14229.4]
  assign _T_12852 = storesToCheck_1_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14230.4]
  assign entriesToCheck_1_9 = _T_12852 & checkBits_1; // @[LoadQueue.scala 141:26:@14231.4]
  assign _T_12854 = storesToCheck_1_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14232.4]
  assign entriesToCheck_1_10 = _T_12854 & checkBits_1; // @[LoadQueue.scala 141:26:@14233.4]
  assign _T_12856 = storesToCheck_1_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14234.4]
  assign entriesToCheck_1_11 = _T_12856 & checkBits_1; // @[LoadQueue.scala 141:26:@14235.4]
  assign _T_12858 = storesToCheck_1_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14236.4]
  assign entriesToCheck_1_12 = _T_12858 & checkBits_1; // @[LoadQueue.scala 141:26:@14237.4]
  assign _T_12860 = storesToCheck_1_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14238.4]
  assign entriesToCheck_1_13 = _T_12860 & checkBits_1; // @[LoadQueue.scala 141:26:@14239.4]
  assign _T_12862 = storesToCheck_1_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14240.4]
  assign entriesToCheck_1_14 = _T_12862 & checkBits_1; // @[LoadQueue.scala 141:26:@14241.4]
  assign _T_12864 = storesToCheck_1_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14242.4]
  assign entriesToCheck_1_15 = _T_12864 & checkBits_1; // @[LoadQueue.scala 141:26:@14243.4]
  assign _T_12866 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14260.4]
  assign entriesToCheck_2_0 = _T_12866 & checkBits_2; // @[LoadQueue.scala 141:26:@14261.4]
  assign _T_12868 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14262.4]
  assign entriesToCheck_2_1 = _T_12868 & checkBits_2; // @[LoadQueue.scala 141:26:@14263.4]
  assign _T_12870 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14264.4]
  assign entriesToCheck_2_2 = _T_12870 & checkBits_2; // @[LoadQueue.scala 141:26:@14265.4]
  assign _T_12872 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14266.4]
  assign entriesToCheck_2_3 = _T_12872 & checkBits_2; // @[LoadQueue.scala 141:26:@14267.4]
  assign _T_12874 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14268.4]
  assign entriesToCheck_2_4 = _T_12874 & checkBits_2; // @[LoadQueue.scala 141:26:@14269.4]
  assign _T_12876 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14270.4]
  assign entriesToCheck_2_5 = _T_12876 & checkBits_2; // @[LoadQueue.scala 141:26:@14271.4]
  assign _T_12878 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14272.4]
  assign entriesToCheck_2_6 = _T_12878 & checkBits_2; // @[LoadQueue.scala 141:26:@14273.4]
  assign _T_12880 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14274.4]
  assign entriesToCheck_2_7 = _T_12880 & checkBits_2; // @[LoadQueue.scala 141:26:@14275.4]
  assign _T_12882 = storesToCheck_2_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14276.4]
  assign entriesToCheck_2_8 = _T_12882 & checkBits_2; // @[LoadQueue.scala 141:26:@14277.4]
  assign _T_12884 = storesToCheck_2_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14278.4]
  assign entriesToCheck_2_9 = _T_12884 & checkBits_2; // @[LoadQueue.scala 141:26:@14279.4]
  assign _T_12886 = storesToCheck_2_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14280.4]
  assign entriesToCheck_2_10 = _T_12886 & checkBits_2; // @[LoadQueue.scala 141:26:@14281.4]
  assign _T_12888 = storesToCheck_2_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14282.4]
  assign entriesToCheck_2_11 = _T_12888 & checkBits_2; // @[LoadQueue.scala 141:26:@14283.4]
  assign _T_12890 = storesToCheck_2_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14284.4]
  assign entriesToCheck_2_12 = _T_12890 & checkBits_2; // @[LoadQueue.scala 141:26:@14285.4]
  assign _T_12892 = storesToCheck_2_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14286.4]
  assign entriesToCheck_2_13 = _T_12892 & checkBits_2; // @[LoadQueue.scala 141:26:@14287.4]
  assign _T_12894 = storesToCheck_2_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14288.4]
  assign entriesToCheck_2_14 = _T_12894 & checkBits_2; // @[LoadQueue.scala 141:26:@14289.4]
  assign _T_12896 = storesToCheck_2_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14290.4]
  assign entriesToCheck_2_15 = _T_12896 & checkBits_2; // @[LoadQueue.scala 141:26:@14291.4]
  assign _T_12898 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14308.4]
  assign entriesToCheck_3_0 = _T_12898 & checkBits_3; // @[LoadQueue.scala 141:26:@14309.4]
  assign _T_12900 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14310.4]
  assign entriesToCheck_3_1 = _T_12900 & checkBits_3; // @[LoadQueue.scala 141:26:@14311.4]
  assign _T_12902 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14312.4]
  assign entriesToCheck_3_2 = _T_12902 & checkBits_3; // @[LoadQueue.scala 141:26:@14313.4]
  assign _T_12904 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14314.4]
  assign entriesToCheck_3_3 = _T_12904 & checkBits_3; // @[LoadQueue.scala 141:26:@14315.4]
  assign _T_12906 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14316.4]
  assign entriesToCheck_3_4 = _T_12906 & checkBits_3; // @[LoadQueue.scala 141:26:@14317.4]
  assign _T_12908 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14318.4]
  assign entriesToCheck_3_5 = _T_12908 & checkBits_3; // @[LoadQueue.scala 141:26:@14319.4]
  assign _T_12910 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14320.4]
  assign entriesToCheck_3_6 = _T_12910 & checkBits_3; // @[LoadQueue.scala 141:26:@14321.4]
  assign _T_12912 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14322.4]
  assign entriesToCheck_3_7 = _T_12912 & checkBits_3; // @[LoadQueue.scala 141:26:@14323.4]
  assign _T_12914 = storesToCheck_3_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14324.4]
  assign entriesToCheck_3_8 = _T_12914 & checkBits_3; // @[LoadQueue.scala 141:26:@14325.4]
  assign _T_12916 = storesToCheck_3_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14326.4]
  assign entriesToCheck_3_9 = _T_12916 & checkBits_3; // @[LoadQueue.scala 141:26:@14327.4]
  assign _T_12918 = storesToCheck_3_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14328.4]
  assign entriesToCheck_3_10 = _T_12918 & checkBits_3; // @[LoadQueue.scala 141:26:@14329.4]
  assign _T_12920 = storesToCheck_3_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14330.4]
  assign entriesToCheck_3_11 = _T_12920 & checkBits_3; // @[LoadQueue.scala 141:26:@14331.4]
  assign _T_12922 = storesToCheck_3_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14332.4]
  assign entriesToCheck_3_12 = _T_12922 & checkBits_3; // @[LoadQueue.scala 141:26:@14333.4]
  assign _T_12924 = storesToCheck_3_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14334.4]
  assign entriesToCheck_3_13 = _T_12924 & checkBits_3; // @[LoadQueue.scala 141:26:@14335.4]
  assign _T_12926 = storesToCheck_3_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14336.4]
  assign entriesToCheck_3_14 = _T_12926 & checkBits_3; // @[LoadQueue.scala 141:26:@14337.4]
  assign _T_12928 = storesToCheck_3_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14338.4]
  assign entriesToCheck_3_15 = _T_12928 & checkBits_3; // @[LoadQueue.scala 141:26:@14339.4]
  assign _T_12930 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14356.4]
  assign entriesToCheck_4_0 = _T_12930 & checkBits_4; // @[LoadQueue.scala 141:26:@14357.4]
  assign _T_12932 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14358.4]
  assign entriesToCheck_4_1 = _T_12932 & checkBits_4; // @[LoadQueue.scala 141:26:@14359.4]
  assign _T_12934 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14360.4]
  assign entriesToCheck_4_2 = _T_12934 & checkBits_4; // @[LoadQueue.scala 141:26:@14361.4]
  assign _T_12936 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14362.4]
  assign entriesToCheck_4_3 = _T_12936 & checkBits_4; // @[LoadQueue.scala 141:26:@14363.4]
  assign _T_12938 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14364.4]
  assign entriesToCheck_4_4 = _T_12938 & checkBits_4; // @[LoadQueue.scala 141:26:@14365.4]
  assign _T_12940 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14366.4]
  assign entriesToCheck_4_5 = _T_12940 & checkBits_4; // @[LoadQueue.scala 141:26:@14367.4]
  assign _T_12942 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14368.4]
  assign entriesToCheck_4_6 = _T_12942 & checkBits_4; // @[LoadQueue.scala 141:26:@14369.4]
  assign _T_12944 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14370.4]
  assign entriesToCheck_4_7 = _T_12944 & checkBits_4; // @[LoadQueue.scala 141:26:@14371.4]
  assign _T_12946 = storesToCheck_4_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14372.4]
  assign entriesToCheck_4_8 = _T_12946 & checkBits_4; // @[LoadQueue.scala 141:26:@14373.4]
  assign _T_12948 = storesToCheck_4_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14374.4]
  assign entriesToCheck_4_9 = _T_12948 & checkBits_4; // @[LoadQueue.scala 141:26:@14375.4]
  assign _T_12950 = storesToCheck_4_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14376.4]
  assign entriesToCheck_4_10 = _T_12950 & checkBits_4; // @[LoadQueue.scala 141:26:@14377.4]
  assign _T_12952 = storesToCheck_4_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14378.4]
  assign entriesToCheck_4_11 = _T_12952 & checkBits_4; // @[LoadQueue.scala 141:26:@14379.4]
  assign _T_12954 = storesToCheck_4_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14380.4]
  assign entriesToCheck_4_12 = _T_12954 & checkBits_4; // @[LoadQueue.scala 141:26:@14381.4]
  assign _T_12956 = storesToCheck_4_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14382.4]
  assign entriesToCheck_4_13 = _T_12956 & checkBits_4; // @[LoadQueue.scala 141:26:@14383.4]
  assign _T_12958 = storesToCheck_4_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14384.4]
  assign entriesToCheck_4_14 = _T_12958 & checkBits_4; // @[LoadQueue.scala 141:26:@14385.4]
  assign _T_12960 = storesToCheck_4_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14386.4]
  assign entriesToCheck_4_15 = _T_12960 & checkBits_4; // @[LoadQueue.scala 141:26:@14387.4]
  assign _T_12962 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14404.4]
  assign entriesToCheck_5_0 = _T_12962 & checkBits_5; // @[LoadQueue.scala 141:26:@14405.4]
  assign _T_12964 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14406.4]
  assign entriesToCheck_5_1 = _T_12964 & checkBits_5; // @[LoadQueue.scala 141:26:@14407.4]
  assign _T_12966 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14408.4]
  assign entriesToCheck_5_2 = _T_12966 & checkBits_5; // @[LoadQueue.scala 141:26:@14409.4]
  assign _T_12968 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14410.4]
  assign entriesToCheck_5_3 = _T_12968 & checkBits_5; // @[LoadQueue.scala 141:26:@14411.4]
  assign _T_12970 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14412.4]
  assign entriesToCheck_5_4 = _T_12970 & checkBits_5; // @[LoadQueue.scala 141:26:@14413.4]
  assign _T_12972 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14414.4]
  assign entriesToCheck_5_5 = _T_12972 & checkBits_5; // @[LoadQueue.scala 141:26:@14415.4]
  assign _T_12974 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14416.4]
  assign entriesToCheck_5_6 = _T_12974 & checkBits_5; // @[LoadQueue.scala 141:26:@14417.4]
  assign _T_12976 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14418.4]
  assign entriesToCheck_5_7 = _T_12976 & checkBits_5; // @[LoadQueue.scala 141:26:@14419.4]
  assign _T_12978 = storesToCheck_5_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14420.4]
  assign entriesToCheck_5_8 = _T_12978 & checkBits_5; // @[LoadQueue.scala 141:26:@14421.4]
  assign _T_12980 = storesToCheck_5_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14422.4]
  assign entriesToCheck_5_9 = _T_12980 & checkBits_5; // @[LoadQueue.scala 141:26:@14423.4]
  assign _T_12982 = storesToCheck_5_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14424.4]
  assign entriesToCheck_5_10 = _T_12982 & checkBits_5; // @[LoadQueue.scala 141:26:@14425.4]
  assign _T_12984 = storesToCheck_5_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14426.4]
  assign entriesToCheck_5_11 = _T_12984 & checkBits_5; // @[LoadQueue.scala 141:26:@14427.4]
  assign _T_12986 = storesToCheck_5_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14428.4]
  assign entriesToCheck_5_12 = _T_12986 & checkBits_5; // @[LoadQueue.scala 141:26:@14429.4]
  assign _T_12988 = storesToCheck_5_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14430.4]
  assign entriesToCheck_5_13 = _T_12988 & checkBits_5; // @[LoadQueue.scala 141:26:@14431.4]
  assign _T_12990 = storesToCheck_5_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14432.4]
  assign entriesToCheck_5_14 = _T_12990 & checkBits_5; // @[LoadQueue.scala 141:26:@14433.4]
  assign _T_12992 = storesToCheck_5_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14434.4]
  assign entriesToCheck_5_15 = _T_12992 & checkBits_5; // @[LoadQueue.scala 141:26:@14435.4]
  assign _T_12994 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14452.4]
  assign entriesToCheck_6_0 = _T_12994 & checkBits_6; // @[LoadQueue.scala 141:26:@14453.4]
  assign _T_12996 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14454.4]
  assign entriesToCheck_6_1 = _T_12996 & checkBits_6; // @[LoadQueue.scala 141:26:@14455.4]
  assign _T_12998 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14456.4]
  assign entriesToCheck_6_2 = _T_12998 & checkBits_6; // @[LoadQueue.scala 141:26:@14457.4]
  assign _T_13000 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14458.4]
  assign entriesToCheck_6_3 = _T_13000 & checkBits_6; // @[LoadQueue.scala 141:26:@14459.4]
  assign _T_13002 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14460.4]
  assign entriesToCheck_6_4 = _T_13002 & checkBits_6; // @[LoadQueue.scala 141:26:@14461.4]
  assign _T_13004 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14462.4]
  assign entriesToCheck_6_5 = _T_13004 & checkBits_6; // @[LoadQueue.scala 141:26:@14463.4]
  assign _T_13006 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14464.4]
  assign entriesToCheck_6_6 = _T_13006 & checkBits_6; // @[LoadQueue.scala 141:26:@14465.4]
  assign _T_13008 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14466.4]
  assign entriesToCheck_6_7 = _T_13008 & checkBits_6; // @[LoadQueue.scala 141:26:@14467.4]
  assign _T_13010 = storesToCheck_6_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14468.4]
  assign entriesToCheck_6_8 = _T_13010 & checkBits_6; // @[LoadQueue.scala 141:26:@14469.4]
  assign _T_13012 = storesToCheck_6_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14470.4]
  assign entriesToCheck_6_9 = _T_13012 & checkBits_6; // @[LoadQueue.scala 141:26:@14471.4]
  assign _T_13014 = storesToCheck_6_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14472.4]
  assign entriesToCheck_6_10 = _T_13014 & checkBits_6; // @[LoadQueue.scala 141:26:@14473.4]
  assign _T_13016 = storesToCheck_6_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14474.4]
  assign entriesToCheck_6_11 = _T_13016 & checkBits_6; // @[LoadQueue.scala 141:26:@14475.4]
  assign _T_13018 = storesToCheck_6_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14476.4]
  assign entriesToCheck_6_12 = _T_13018 & checkBits_6; // @[LoadQueue.scala 141:26:@14477.4]
  assign _T_13020 = storesToCheck_6_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14478.4]
  assign entriesToCheck_6_13 = _T_13020 & checkBits_6; // @[LoadQueue.scala 141:26:@14479.4]
  assign _T_13022 = storesToCheck_6_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14480.4]
  assign entriesToCheck_6_14 = _T_13022 & checkBits_6; // @[LoadQueue.scala 141:26:@14481.4]
  assign _T_13024 = storesToCheck_6_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14482.4]
  assign entriesToCheck_6_15 = _T_13024 & checkBits_6; // @[LoadQueue.scala 141:26:@14483.4]
  assign _T_13026 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14500.4]
  assign entriesToCheck_7_0 = _T_13026 & checkBits_7; // @[LoadQueue.scala 141:26:@14501.4]
  assign _T_13028 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14502.4]
  assign entriesToCheck_7_1 = _T_13028 & checkBits_7; // @[LoadQueue.scala 141:26:@14503.4]
  assign _T_13030 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14504.4]
  assign entriesToCheck_7_2 = _T_13030 & checkBits_7; // @[LoadQueue.scala 141:26:@14505.4]
  assign _T_13032 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14506.4]
  assign entriesToCheck_7_3 = _T_13032 & checkBits_7; // @[LoadQueue.scala 141:26:@14507.4]
  assign _T_13034 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14508.4]
  assign entriesToCheck_7_4 = _T_13034 & checkBits_7; // @[LoadQueue.scala 141:26:@14509.4]
  assign _T_13036 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14510.4]
  assign entriesToCheck_7_5 = _T_13036 & checkBits_7; // @[LoadQueue.scala 141:26:@14511.4]
  assign _T_13038 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14512.4]
  assign entriesToCheck_7_6 = _T_13038 & checkBits_7; // @[LoadQueue.scala 141:26:@14513.4]
  assign _T_13040 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14514.4]
  assign entriesToCheck_7_7 = _T_13040 & checkBits_7; // @[LoadQueue.scala 141:26:@14515.4]
  assign _T_13042 = storesToCheck_7_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14516.4]
  assign entriesToCheck_7_8 = _T_13042 & checkBits_7; // @[LoadQueue.scala 141:26:@14517.4]
  assign _T_13044 = storesToCheck_7_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14518.4]
  assign entriesToCheck_7_9 = _T_13044 & checkBits_7; // @[LoadQueue.scala 141:26:@14519.4]
  assign _T_13046 = storesToCheck_7_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14520.4]
  assign entriesToCheck_7_10 = _T_13046 & checkBits_7; // @[LoadQueue.scala 141:26:@14521.4]
  assign _T_13048 = storesToCheck_7_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14522.4]
  assign entriesToCheck_7_11 = _T_13048 & checkBits_7; // @[LoadQueue.scala 141:26:@14523.4]
  assign _T_13050 = storesToCheck_7_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14524.4]
  assign entriesToCheck_7_12 = _T_13050 & checkBits_7; // @[LoadQueue.scala 141:26:@14525.4]
  assign _T_13052 = storesToCheck_7_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14526.4]
  assign entriesToCheck_7_13 = _T_13052 & checkBits_7; // @[LoadQueue.scala 141:26:@14527.4]
  assign _T_13054 = storesToCheck_7_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14528.4]
  assign entriesToCheck_7_14 = _T_13054 & checkBits_7; // @[LoadQueue.scala 141:26:@14529.4]
  assign _T_13056 = storesToCheck_7_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14530.4]
  assign entriesToCheck_7_15 = _T_13056 & checkBits_7; // @[LoadQueue.scala 141:26:@14531.4]
  assign _T_13058 = storesToCheck_8_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14548.4]
  assign entriesToCheck_8_0 = _T_13058 & checkBits_8; // @[LoadQueue.scala 141:26:@14549.4]
  assign _T_13060 = storesToCheck_8_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14550.4]
  assign entriesToCheck_8_1 = _T_13060 & checkBits_8; // @[LoadQueue.scala 141:26:@14551.4]
  assign _T_13062 = storesToCheck_8_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14552.4]
  assign entriesToCheck_8_2 = _T_13062 & checkBits_8; // @[LoadQueue.scala 141:26:@14553.4]
  assign _T_13064 = storesToCheck_8_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14554.4]
  assign entriesToCheck_8_3 = _T_13064 & checkBits_8; // @[LoadQueue.scala 141:26:@14555.4]
  assign _T_13066 = storesToCheck_8_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14556.4]
  assign entriesToCheck_8_4 = _T_13066 & checkBits_8; // @[LoadQueue.scala 141:26:@14557.4]
  assign _T_13068 = storesToCheck_8_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14558.4]
  assign entriesToCheck_8_5 = _T_13068 & checkBits_8; // @[LoadQueue.scala 141:26:@14559.4]
  assign _T_13070 = storesToCheck_8_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14560.4]
  assign entriesToCheck_8_6 = _T_13070 & checkBits_8; // @[LoadQueue.scala 141:26:@14561.4]
  assign _T_13072 = storesToCheck_8_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14562.4]
  assign entriesToCheck_8_7 = _T_13072 & checkBits_8; // @[LoadQueue.scala 141:26:@14563.4]
  assign _T_13074 = storesToCheck_8_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14564.4]
  assign entriesToCheck_8_8 = _T_13074 & checkBits_8; // @[LoadQueue.scala 141:26:@14565.4]
  assign _T_13076 = storesToCheck_8_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14566.4]
  assign entriesToCheck_8_9 = _T_13076 & checkBits_8; // @[LoadQueue.scala 141:26:@14567.4]
  assign _T_13078 = storesToCheck_8_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14568.4]
  assign entriesToCheck_8_10 = _T_13078 & checkBits_8; // @[LoadQueue.scala 141:26:@14569.4]
  assign _T_13080 = storesToCheck_8_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14570.4]
  assign entriesToCheck_8_11 = _T_13080 & checkBits_8; // @[LoadQueue.scala 141:26:@14571.4]
  assign _T_13082 = storesToCheck_8_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14572.4]
  assign entriesToCheck_8_12 = _T_13082 & checkBits_8; // @[LoadQueue.scala 141:26:@14573.4]
  assign _T_13084 = storesToCheck_8_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14574.4]
  assign entriesToCheck_8_13 = _T_13084 & checkBits_8; // @[LoadQueue.scala 141:26:@14575.4]
  assign _T_13086 = storesToCheck_8_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14576.4]
  assign entriesToCheck_8_14 = _T_13086 & checkBits_8; // @[LoadQueue.scala 141:26:@14577.4]
  assign _T_13088 = storesToCheck_8_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14578.4]
  assign entriesToCheck_8_15 = _T_13088 & checkBits_8; // @[LoadQueue.scala 141:26:@14579.4]
  assign _T_13090 = storesToCheck_9_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14596.4]
  assign entriesToCheck_9_0 = _T_13090 & checkBits_9; // @[LoadQueue.scala 141:26:@14597.4]
  assign _T_13092 = storesToCheck_9_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14598.4]
  assign entriesToCheck_9_1 = _T_13092 & checkBits_9; // @[LoadQueue.scala 141:26:@14599.4]
  assign _T_13094 = storesToCheck_9_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14600.4]
  assign entriesToCheck_9_2 = _T_13094 & checkBits_9; // @[LoadQueue.scala 141:26:@14601.4]
  assign _T_13096 = storesToCheck_9_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14602.4]
  assign entriesToCheck_9_3 = _T_13096 & checkBits_9; // @[LoadQueue.scala 141:26:@14603.4]
  assign _T_13098 = storesToCheck_9_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14604.4]
  assign entriesToCheck_9_4 = _T_13098 & checkBits_9; // @[LoadQueue.scala 141:26:@14605.4]
  assign _T_13100 = storesToCheck_9_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14606.4]
  assign entriesToCheck_9_5 = _T_13100 & checkBits_9; // @[LoadQueue.scala 141:26:@14607.4]
  assign _T_13102 = storesToCheck_9_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14608.4]
  assign entriesToCheck_9_6 = _T_13102 & checkBits_9; // @[LoadQueue.scala 141:26:@14609.4]
  assign _T_13104 = storesToCheck_9_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14610.4]
  assign entriesToCheck_9_7 = _T_13104 & checkBits_9; // @[LoadQueue.scala 141:26:@14611.4]
  assign _T_13106 = storesToCheck_9_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14612.4]
  assign entriesToCheck_9_8 = _T_13106 & checkBits_9; // @[LoadQueue.scala 141:26:@14613.4]
  assign _T_13108 = storesToCheck_9_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14614.4]
  assign entriesToCheck_9_9 = _T_13108 & checkBits_9; // @[LoadQueue.scala 141:26:@14615.4]
  assign _T_13110 = storesToCheck_9_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14616.4]
  assign entriesToCheck_9_10 = _T_13110 & checkBits_9; // @[LoadQueue.scala 141:26:@14617.4]
  assign _T_13112 = storesToCheck_9_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14618.4]
  assign entriesToCheck_9_11 = _T_13112 & checkBits_9; // @[LoadQueue.scala 141:26:@14619.4]
  assign _T_13114 = storesToCheck_9_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14620.4]
  assign entriesToCheck_9_12 = _T_13114 & checkBits_9; // @[LoadQueue.scala 141:26:@14621.4]
  assign _T_13116 = storesToCheck_9_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14622.4]
  assign entriesToCheck_9_13 = _T_13116 & checkBits_9; // @[LoadQueue.scala 141:26:@14623.4]
  assign _T_13118 = storesToCheck_9_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14624.4]
  assign entriesToCheck_9_14 = _T_13118 & checkBits_9; // @[LoadQueue.scala 141:26:@14625.4]
  assign _T_13120 = storesToCheck_9_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14626.4]
  assign entriesToCheck_9_15 = _T_13120 & checkBits_9; // @[LoadQueue.scala 141:26:@14627.4]
  assign _T_13122 = storesToCheck_10_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14644.4]
  assign entriesToCheck_10_0 = _T_13122 & checkBits_10; // @[LoadQueue.scala 141:26:@14645.4]
  assign _T_13124 = storesToCheck_10_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14646.4]
  assign entriesToCheck_10_1 = _T_13124 & checkBits_10; // @[LoadQueue.scala 141:26:@14647.4]
  assign _T_13126 = storesToCheck_10_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14648.4]
  assign entriesToCheck_10_2 = _T_13126 & checkBits_10; // @[LoadQueue.scala 141:26:@14649.4]
  assign _T_13128 = storesToCheck_10_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14650.4]
  assign entriesToCheck_10_3 = _T_13128 & checkBits_10; // @[LoadQueue.scala 141:26:@14651.4]
  assign _T_13130 = storesToCheck_10_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14652.4]
  assign entriesToCheck_10_4 = _T_13130 & checkBits_10; // @[LoadQueue.scala 141:26:@14653.4]
  assign _T_13132 = storesToCheck_10_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14654.4]
  assign entriesToCheck_10_5 = _T_13132 & checkBits_10; // @[LoadQueue.scala 141:26:@14655.4]
  assign _T_13134 = storesToCheck_10_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14656.4]
  assign entriesToCheck_10_6 = _T_13134 & checkBits_10; // @[LoadQueue.scala 141:26:@14657.4]
  assign _T_13136 = storesToCheck_10_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14658.4]
  assign entriesToCheck_10_7 = _T_13136 & checkBits_10; // @[LoadQueue.scala 141:26:@14659.4]
  assign _T_13138 = storesToCheck_10_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14660.4]
  assign entriesToCheck_10_8 = _T_13138 & checkBits_10; // @[LoadQueue.scala 141:26:@14661.4]
  assign _T_13140 = storesToCheck_10_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14662.4]
  assign entriesToCheck_10_9 = _T_13140 & checkBits_10; // @[LoadQueue.scala 141:26:@14663.4]
  assign _T_13142 = storesToCheck_10_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14664.4]
  assign entriesToCheck_10_10 = _T_13142 & checkBits_10; // @[LoadQueue.scala 141:26:@14665.4]
  assign _T_13144 = storesToCheck_10_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14666.4]
  assign entriesToCheck_10_11 = _T_13144 & checkBits_10; // @[LoadQueue.scala 141:26:@14667.4]
  assign _T_13146 = storesToCheck_10_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14668.4]
  assign entriesToCheck_10_12 = _T_13146 & checkBits_10; // @[LoadQueue.scala 141:26:@14669.4]
  assign _T_13148 = storesToCheck_10_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14670.4]
  assign entriesToCheck_10_13 = _T_13148 & checkBits_10; // @[LoadQueue.scala 141:26:@14671.4]
  assign _T_13150 = storesToCheck_10_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14672.4]
  assign entriesToCheck_10_14 = _T_13150 & checkBits_10; // @[LoadQueue.scala 141:26:@14673.4]
  assign _T_13152 = storesToCheck_10_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14674.4]
  assign entriesToCheck_10_15 = _T_13152 & checkBits_10; // @[LoadQueue.scala 141:26:@14675.4]
  assign _T_13154 = storesToCheck_11_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14692.4]
  assign entriesToCheck_11_0 = _T_13154 & checkBits_11; // @[LoadQueue.scala 141:26:@14693.4]
  assign _T_13156 = storesToCheck_11_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14694.4]
  assign entriesToCheck_11_1 = _T_13156 & checkBits_11; // @[LoadQueue.scala 141:26:@14695.4]
  assign _T_13158 = storesToCheck_11_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14696.4]
  assign entriesToCheck_11_2 = _T_13158 & checkBits_11; // @[LoadQueue.scala 141:26:@14697.4]
  assign _T_13160 = storesToCheck_11_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14698.4]
  assign entriesToCheck_11_3 = _T_13160 & checkBits_11; // @[LoadQueue.scala 141:26:@14699.4]
  assign _T_13162 = storesToCheck_11_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14700.4]
  assign entriesToCheck_11_4 = _T_13162 & checkBits_11; // @[LoadQueue.scala 141:26:@14701.4]
  assign _T_13164 = storesToCheck_11_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14702.4]
  assign entriesToCheck_11_5 = _T_13164 & checkBits_11; // @[LoadQueue.scala 141:26:@14703.4]
  assign _T_13166 = storesToCheck_11_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14704.4]
  assign entriesToCheck_11_6 = _T_13166 & checkBits_11; // @[LoadQueue.scala 141:26:@14705.4]
  assign _T_13168 = storesToCheck_11_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14706.4]
  assign entriesToCheck_11_7 = _T_13168 & checkBits_11; // @[LoadQueue.scala 141:26:@14707.4]
  assign _T_13170 = storesToCheck_11_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14708.4]
  assign entriesToCheck_11_8 = _T_13170 & checkBits_11; // @[LoadQueue.scala 141:26:@14709.4]
  assign _T_13172 = storesToCheck_11_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14710.4]
  assign entriesToCheck_11_9 = _T_13172 & checkBits_11; // @[LoadQueue.scala 141:26:@14711.4]
  assign _T_13174 = storesToCheck_11_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14712.4]
  assign entriesToCheck_11_10 = _T_13174 & checkBits_11; // @[LoadQueue.scala 141:26:@14713.4]
  assign _T_13176 = storesToCheck_11_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14714.4]
  assign entriesToCheck_11_11 = _T_13176 & checkBits_11; // @[LoadQueue.scala 141:26:@14715.4]
  assign _T_13178 = storesToCheck_11_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14716.4]
  assign entriesToCheck_11_12 = _T_13178 & checkBits_11; // @[LoadQueue.scala 141:26:@14717.4]
  assign _T_13180 = storesToCheck_11_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14718.4]
  assign entriesToCheck_11_13 = _T_13180 & checkBits_11; // @[LoadQueue.scala 141:26:@14719.4]
  assign _T_13182 = storesToCheck_11_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14720.4]
  assign entriesToCheck_11_14 = _T_13182 & checkBits_11; // @[LoadQueue.scala 141:26:@14721.4]
  assign _T_13184 = storesToCheck_11_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14722.4]
  assign entriesToCheck_11_15 = _T_13184 & checkBits_11; // @[LoadQueue.scala 141:26:@14723.4]
  assign _T_13186 = storesToCheck_12_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14740.4]
  assign entriesToCheck_12_0 = _T_13186 & checkBits_12; // @[LoadQueue.scala 141:26:@14741.4]
  assign _T_13188 = storesToCheck_12_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14742.4]
  assign entriesToCheck_12_1 = _T_13188 & checkBits_12; // @[LoadQueue.scala 141:26:@14743.4]
  assign _T_13190 = storesToCheck_12_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14744.4]
  assign entriesToCheck_12_2 = _T_13190 & checkBits_12; // @[LoadQueue.scala 141:26:@14745.4]
  assign _T_13192 = storesToCheck_12_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14746.4]
  assign entriesToCheck_12_3 = _T_13192 & checkBits_12; // @[LoadQueue.scala 141:26:@14747.4]
  assign _T_13194 = storesToCheck_12_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14748.4]
  assign entriesToCheck_12_4 = _T_13194 & checkBits_12; // @[LoadQueue.scala 141:26:@14749.4]
  assign _T_13196 = storesToCheck_12_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14750.4]
  assign entriesToCheck_12_5 = _T_13196 & checkBits_12; // @[LoadQueue.scala 141:26:@14751.4]
  assign _T_13198 = storesToCheck_12_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14752.4]
  assign entriesToCheck_12_6 = _T_13198 & checkBits_12; // @[LoadQueue.scala 141:26:@14753.4]
  assign _T_13200 = storesToCheck_12_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14754.4]
  assign entriesToCheck_12_7 = _T_13200 & checkBits_12; // @[LoadQueue.scala 141:26:@14755.4]
  assign _T_13202 = storesToCheck_12_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14756.4]
  assign entriesToCheck_12_8 = _T_13202 & checkBits_12; // @[LoadQueue.scala 141:26:@14757.4]
  assign _T_13204 = storesToCheck_12_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14758.4]
  assign entriesToCheck_12_9 = _T_13204 & checkBits_12; // @[LoadQueue.scala 141:26:@14759.4]
  assign _T_13206 = storesToCheck_12_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14760.4]
  assign entriesToCheck_12_10 = _T_13206 & checkBits_12; // @[LoadQueue.scala 141:26:@14761.4]
  assign _T_13208 = storesToCheck_12_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14762.4]
  assign entriesToCheck_12_11 = _T_13208 & checkBits_12; // @[LoadQueue.scala 141:26:@14763.4]
  assign _T_13210 = storesToCheck_12_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14764.4]
  assign entriesToCheck_12_12 = _T_13210 & checkBits_12; // @[LoadQueue.scala 141:26:@14765.4]
  assign _T_13212 = storesToCheck_12_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14766.4]
  assign entriesToCheck_12_13 = _T_13212 & checkBits_12; // @[LoadQueue.scala 141:26:@14767.4]
  assign _T_13214 = storesToCheck_12_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14768.4]
  assign entriesToCheck_12_14 = _T_13214 & checkBits_12; // @[LoadQueue.scala 141:26:@14769.4]
  assign _T_13216 = storesToCheck_12_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14770.4]
  assign entriesToCheck_12_15 = _T_13216 & checkBits_12; // @[LoadQueue.scala 141:26:@14771.4]
  assign _T_13218 = storesToCheck_13_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14788.4]
  assign entriesToCheck_13_0 = _T_13218 & checkBits_13; // @[LoadQueue.scala 141:26:@14789.4]
  assign _T_13220 = storesToCheck_13_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14790.4]
  assign entriesToCheck_13_1 = _T_13220 & checkBits_13; // @[LoadQueue.scala 141:26:@14791.4]
  assign _T_13222 = storesToCheck_13_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14792.4]
  assign entriesToCheck_13_2 = _T_13222 & checkBits_13; // @[LoadQueue.scala 141:26:@14793.4]
  assign _T_13224 = storesToCheck_13_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14794.4]
  assign entriesToCheck_13_3 = _T_13224 & checkBits_13; // @[LoadQueue.scala 141:26:@14795.4]
  assign _T_13226 = storesToCheck_13_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14796.4]
  assign entriesToCheck_13_4 = _T_13226 & checkBits_13; // @[LoadQueue.scala 141:26:@14797.4]
  assign _T_13228 = storesToCheck_13_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14798.4]
  assign entriesToCheck_13_5 = _T_13228 & checkBits_13; // @[LoadQueue.scala 141:26:@14799.4]
  assign _T_13230 = storesToCheck_13_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14800.4]
  assign entriesToCheck_13_6 = _T_13230 & checkBits_13; // @[LoadQueue.scala 141:26:@14801.4]
  assign _T_13232 = storesToCheck_13_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14802.4]
  assign entriesToCheck_13_7 = _T_13232 & checkBits_13; // @[LoadQueue.scala 141:26:@14803.4]
  assign _T_13234 = storesToCheck_13_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14804.4]
  assign entriesToCheck_13_8 = _T_13234 & checkBits_13; // @[LoadQueue.scala 141:26:@14805.4]
  assign _T_13236 = storesToCheck_13_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14806.4]
  assign entriesToCheck_13_9 = _T_13236 & checkBits_13; // @[LoadQueue.scala 141:26:@14807.4]
  assign _T_13238 = storesToCheck_13_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14808.4]
  assign entriesToCheck_13_10 = _T_13238 & checkBits_13; // @[LoadQueue.scala 141:26:@14809.4]
  assign _T_13240 = storesToCheck_13_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14810.4]
  assign entriesToCheck_13_11 = _T_13240 & checkBits_13; // @[LoadQueue.scala 141:26:@14811.4]
  assign _T_13242 = storesToCheck_13_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14812.4]
  assign entriesToCheck_13_12 = _T_13242 & checkBits_13; // @[LoadQueue.scala 141:26:@14813.4]
  assign _T_13244 = storesToCheck_13_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14814.4]
  assign entriesToCheck_13_13 = _T_13244 & checkBits_13; // @[LoadQueue.scala 141:26:@14815.4]
  assign _T_13246 = storesToCheck_13_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14816.4]
  assign entriesToCheck_13_14 = _T_13246 & checkBits_13; // @[LoadQueue.scala 141:26:@14817.4]
  assign _T_13248 = storesToCheck_13_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14818.4]
  assign entriesToCheck_13_15 = _T_13248 & checkBits_13; // @[LoadQueue.scala 141:26:@14819.4]
  assign _T_13250 = storesToCheck_14_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14836.4]
  assign entriesToCheck_14_0 = _T_13250 & checkBits_14; // @[LoadQueue.scala 141:26:@14837.4]
  assign _T_13252 = storesToCheck_14_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14838.4]
  assign entriesToCheck_14_1 = _T_13252 & checkBits_14; // @[LoadQueue.scala 141:26:@14839.4]
  assign _T_13254 = storesToCheck_14_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14840.4]
  assign entriesToCheck_14_2 = _T_13254 & checkBits_14; // @[LoadQueue.scala 141:26:@14841.4]
  assign _T_13256 = storesToCheck_14_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14842.4]
  assign entriesToCheck_14_3 = _T_13256 & checkBits_14; // @[LoadQueue.scala 141:26:@14843.4]
  assign _T_13258 = storesToCheck_14_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14844.4]
  assign entriesToCheck_14_4 = _T_13258 & checkBits_14; // @[LoadQueue.scala 141:26:@14845.4]
  assign _T_13260 = storesToCheck_14_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14846.4]
  assign entriesToCheck_14_5 = _T_13260 & checkBits_14; // @[LoadQueue.scala 141:26:@14847.4]
  assign _T_13262 = storesToCheck_14_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14848.4]
  assign entriesToCheck_14_6 = _T_13262 & checkBits_14; // @[LoadQueue.scala 141:26:@14849.4]
  assign _T_13264 = storesToCheck_14_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14850.4]
  assign entriesToCheck_14_7 = _T_13264 & checkBits_14; // @[LoadQueue.scala 141:26:@14851.4]
  assign _T_13266 = storesToCheck_14_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14852.4]
  assign entriesToCheck_14_8 = _T_13266 & checkBits_14; // @[LoadQueue.scala 141:26:@14853.4]
  assign _T_13268 = storesToCheck_14_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14854.4]
  assign entriesToCheck_14_9 = _T_13268 & checkBits_14; // @[LoadQueue.scala 141:26:@14855.4]
  assign _T_13270 = storesToCheck_14_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14856.4]
  assign entriesToCheck_14_10 = _T_13270 & checkBits_14; // @[LoadQueue.scala 141:26:@14857.4]
  assign _T_13272 = storesToCheck_14_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14858.4]
  assign entriesToCheck_14_11 = _T_13272 & checkBits_14; // @[LoadQueue.scala 141:26:@14859.4]
  assign _T_13274 = storesToCheck_14_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14860.4]
  assign entriesToCheck_14_12 = _T_13274 & checkBits_14; // @[LoadQueue.scala 141:26:@14861.4]
  assign _T_13276 = storesToCheck_14_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14862.4]
  assign entriesToCheck_14_13 = _T_13276 & checkBits_14; // @[LoadQueue.scala 141:26:@14863.4]
  assign _T_13278 = storesToCheck_14_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14864.4]
  assign entriesToCheck_14_14 = _T_13278 & checkBits_14; // @[LoadQueue.scala 141:26:@14865.4]
  assign _T_13280 = storesToCheck_14_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14866.4]
  assign entriesToCheck_14_15 = _T_13280 & checkBits_14; // @[LoadQueue.scala 141:26:@14867.4]
  assign _T_13282 = storesToCheck_15_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@14884.4]
  assign entriesToCheck_15_0 = _T_13282 & checkBits_15; // @[LoadQueue.scala 141:26:@14885.4]
  assign _T_13284 = storesToCheck_15_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@14886.4]
  assign entriesToCheck_15_1 = _T_13284 & checkBits_15; // @[LoadQueue.scala 141:26:@14887.4]
  assign _T_13286 = storesToCheck_15_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@14888.4]
  assign entriesToCheck_15_2 = _T_13286 & checkBits_15; // @[LoadQueue.scala 141:26:@14889.4]
  assign _T_13288 = storesToCheck_15_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@14890.4]
  assign entriesToCheck_15_3 = _T_13288 & checkBits_15; // @[LoadQueue.scala 141:26:@14891.4]
  assign _T_13290 = storesToCheck_15_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@14892.4]
  assign entriesToCheck_15_4 = _T_13290 & checkBits_15; // @[LoadQueue.scala 141:26:@14893.4]
  assign _T_13292 = storesToCheck_15_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@14894.4]
  assign entriesToCheck_15_5 = _T_13292 & checkBits_15; // @[LoadQueue.scala 141:26:@14895.4]
  assign _T_13294 = storesToCheck_15_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@14896.4]
  assign entriesToCheck_15_6 = _T_13294 & checkBits_15; // @[LoadQueue.scala 141:26:@14897.4]
  assign _T_13296 = storesToCheck_15_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@14898.4]
  assign entriesToCheck_15_7 = _T_13296 & checkBits_15; // @[LoadQueue.scala 141:26:@14899.4]
  assign _T_13298 = storesToCheck_15_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@14900.4]
  assign entriesToCheck_15_8 = _T_13298 & checkBits_15; // @[LoadQueue.scala 141:26:@14901.4]
  assign _T_13300 = storesToCheck_15_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@14902.4]
  assign entriesToCheck_15_9 = _T_13300 & checkBits_15; // @[LoadQueue.scala 141:26:@14903.4]
  assign _T_13302 = storesToCheck_15_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@14904.4]
  assign entriesToCheck_15_10 = _T_13302 & checkBits_15; // @[LoadQueue.scala 141:26:@14905.4]
  assign _T_13304 = storesToCheck_15_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@14906.4]
  assign entriesToCheck_15_11 = _T_13304 & checkBits_15; // @[LoadQueue.scala 141:26:@14907.4]
  assign _T_13306 = storesToCheck_15_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@14908.4]
  assign entriesToCheck_15_12 = _T_13306 & checkBits_15; // @[LoadQueue.scala 141:26:@14909.4]
  assign _T_13308 = storesToCheck_15_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@14910.4]
  assign entriesToCheck_15_13 = _T_13308 & checkBits_15; // @[LoadQueue.scala 141:26:@14911.4]
  assign _T_13310 = storesToCheck_15_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@14912.4]
  assign entriesToCheck_15_14 = _T_13310 & checkBits_15; // @[LoadQueue.scala 141:26:@14913.4]
  assign _T_13312 = storesToCheck_15_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@14914.4]
  assign entriesToCheck_15_15 = _T_13312 & checkBits_15; // @[LoadQueue.scala 141:26:@14915.4]
  assign _T_14544 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@14933.4]
  assign _T_14545 = _T_14544 & addrKnown_0; // @[LoadQueue.scala 152:41:@14934.4]
  assign _T_14546 = addrQ_0 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@14935.4]
  assign conflict_0_0 = _T_14545 & _T_14546; // @[LoadQueue.scala 152:68:@14936.4]
  assign _T_14548 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@14938.4]
  assign _T_14549 = _T_14548 & addrKnown_0; // @[LoadQueue.scala 152:41:@14939.4]
  assign _T_14550 = addrQ_0 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@14940.4]
  assign conflict_0_1 = _T_14549 & _T_14550; // @[LoadQueue.scala 152:68:@14941.4]
  assign _T_14552 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@14943.4]
  assign _T_14553 = _T_14552 & addrKnown_0; // @[LoadQueue.scala 152:41:@14944.4]
  assign _T_14554 = addrQ_0 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@14945.4]
  assign conflict_0_2 = _T_14553 & _T_14554; // @[LoadQueue.scala 152:68:@14946.4]
  assign _T_14556 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@14948.4]
  assign _T_14557 = _T_14556 & addrKnown_0; // @[LoadQueue.scala 152:41:@14949.4]
  assign _T_14558 = addrQ_0 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@14950.4]
  assign conflict_0_3 = _T_14557 & _T_14558; // @[LoadQueue.scala 152:68:@14951.4]
  assign _T_14560 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@14953.4]
  assign _T_14561 = _T_14560 & addrKnown_0; // @[LoadQueue.scala 152:41:@14954.4]
  assign _T_14562 = addrQ_0 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@14955.4]
  assign conflict_0_4 = _T_14561 & _T_14562; // @[LoadQueue.scala 152:68:@14956.4]
  assign _T_14564 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@14958.4]
  assign _T_14565 = _T_14564 & addrKnown_0; // @[LoadQueue.scala 152:41:@14959.4]
  assign _T_14566 = addrQ_0 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@14960.4]
  assign conflict_0_5 = _T_14565 & _T_14566; // @[LoadQueue.scala 152:68:@14961.4]
  assign _T_14568 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@14963.4]
  assign _T_14569 = _T_14568 & addrKnown_0; // @[LoadQueue.scala 152:41:@14964.4]
  assign _T_14570 = addrQ_0 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@14965.4]
  assign conflict_0_6 = _T_14569 & _T_14570; // @[LoadQueue.scala 152:68:@14966.4]
  assign _T_14572 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@14968.4]
  assign _T_14573 = _T_14572 & addrKnown_0; // @[LoadQueue.scala 152:41:@14969.4]
  assign _T_14574 = addrQ_0 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@14970.4]
  assign conflict_0_7 = _T_14573 & _T_14574; // @[LoadQueue.scala 152:68:@14971.4]
  assign _T_14576 = entriesToCheck_0_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@14973.4]
  assign _T_14577 = _T_14576 & addrKnown_0; // @[LoadQueue.scala 152:41:@14974.4]
  assign _T_14578 = addrQ_0 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@14975.4]
  assign conflict_0_8 = _T_14577 & _T_14578; // @[LoadQueue.scala 152:68:@14976.4]
  assign _T_14580 = entriesToCheck_0_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@14978.4]
  assign _T_14581 = _T_14580 & addrKnown_0; // @[LoadQueue.scala 152:41:@14979.4]
  assign _T_14582 = addrQ_0 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@14980.4]
  assign conflict_0_9 = _T_14581 & _T_14582; // @[LoadQueue.scala 152:68:@14981.4]
  assign _T_14584 = entriesToCheck_0_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@14983.4]
  assign _T_14585 = _T_14584 & addrKnown_0; // @[LoadQueue.scala 152:41:@14984.4]
  assign _T_14586 = addrQ_0 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@14985.4]
  assign conflict_0_10 = _T_14585 & _T_14586; // @[LoadQueue.scala 152:68:@14986.4]
  assign _T_14588 = entriesToCheck_0_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@14988.4]
  assign _T_14589 = _T_14588 & addrKnown_0; // @[LoadQueue.scala 152:41:@14989.4]
  assign _T_14590 = addrQ_0 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@14990.4]
  assign conflict_0_11 = _T_14589 & _T_14590; // @[LoadQueue.scala 152:68:@14991.4]
  assign _T_14592 = entriesToCheck_0_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@14993.4]
  assign _T_14593 = _T_14592 & addrKnown_0; // @[LoadQueue.scala 152:41:@14994.4]
  assign _T_14594 = addrQ_0 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@14995.4]
  assign conflict_0_12 = _T_14593 & _T_14594; // @[LoadQueue.scala 152:68:@14996.4]
  assign _T_14596 = entriesToCheck_0_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@14998.4]
  assign _T_14597 = _T_14596 & addrKnown_0; // @[LoadQueue.scala 152:41:@14999.4]
  assign _T_14598 = addrQ_0 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15000.4]
  assign conflict_0_13 = _T_14597 & _T_14598; // @[LoadQueue.scala 152:68:@15001.4]
  assign _T_14600 = entriesToCheck_0_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15003.4]
  assign _T_14601 = _T_14600 & addrKnown_0; // @[LoadQueue.scala 152:41:@15004.4]
  assign _T_14602 = addrQ_0 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15005.4]
  assign conflict_0_14 = _T_14601 & _T_14602; // @[LoadQueue.scala 152:68:@15006.4]
  assign _T_14604 = entriesToCheck_0_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15008.4]
  assign _T_14605 = _T_14604 & addrKnown_0; // @[LoadQueue.scala 152:41:@15009.4]
  assign _T_14606 = addrQ_0 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15010.4]
  assign conflict_0_15 = _T_14605 & _T_14606; // @[LoadQueue.scala 152:68:@15011.4]
  assign _T_14608 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15013.4]
  assign _T_14609 = _T_14608 & addrKnown_1; // @[LoadQueue.scala 152:41:@15014.4]
  assign _T_14610 = addrQ_1 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15015.4]
  assign conflict_1_0 = _T_14609 & _T_14610; // @[LoadQueue.scala 152:68:@15016.4]
  assign _T_14612 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15018.4]
  assign _T_14613 = _T_14612 & addrKnown_1; // @[LoadQueue.scala 152:41:@15019.4]
  assign _T_14614 = addrQ_1 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15020.4]
  assign conflict_1_1 = _T_14613 & _T_14614; // @[LoadQueue.scala 152:68:@15021.4]
  assign _T_14616 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15023.4]
  assign _T_14617 = _T_14616 & addrKnown_1; // @[LoadQueue.scala 152:41:@15024.4]
  assign _T_14618 = addrQ_1 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15025.4]
  assign conflict_1_2 = _T_14617 & _T_14618; // @[LoadQueue.scala 152:68:@15026.4]
  assign _T_14620 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15028.4]
  assign _T_14621 = _T_14620 & addrKnown_1; // @[LoadQueue.scala 152:41:@15029.4]
  assign _T_14622 = addrQ_1 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15030.4]
  assign conflict_1_3 = _T_14621 & _T_14622; // @[LoadQueue.scala 152:68:@15031.4]
  assign _T_14624 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15033.4]
  assign _T_14625 = _T_14624 & addrKnown_1; // @[LoadQueue.scala 152:41:@15034.4]
  assign _T_14626 = addrQ_1 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15035.4]
  assign conflict_1_4 = _T_14625 & _T_14626; // @[LoadQueue.scala 152:68:@15036.4]
  assign _T_14628 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15038.4]
  assign _T_14629 = _T_14628 & addrKnown_1; // @[LoadQueue.scala 152:41:@15039.4]
  assign _T_14630 = addrQ_1 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15040.4]
  assign conflict_1_5 = _T_14629 & _T_14630; // @[LoadQueue.scala 152:68:@15041.4]
  assign _T_14632 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15043.4]
  assign _T_14633 = _T_14632 & addrKnown_1; // @[LoadQueue.scala 152:41:@15044.4]
  assign _T_14634 = addrQ_1 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15045.4]
  assign conflict_1_6 = _T_14633 & _T_14634; // @[LoadQueue.scala 152:68:@15046.4]
  assign _T_14636 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15048.4]
  assign _T_14637 = _T_14636 & addrKnown_1; // @[LoadQueue.scala 152:41:@15049.4]
  assign _T_14638 = addrQ_1 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15050.4]
  assign conflict_1_7 = _T_14637 & _T_14638; // @[LoadQueue.scala 152:68:@15051.4]
  assign _T_14640 = entriesToCheck_1_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15053.4]
  assign _T_14641 = _T_14640 & addrKnown_1; // @[LoadQueue.scala 152:41:@15054.4]
  assign _T_14642 = addrQ_1 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15055.4]
  assign conflict_1_8 = _T_14641 & _T_14642; // @[LoadQueue.scala 152:68:@15056.4]
  assign _T_14644 = entriesToCheck_1_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15058.4]
  assign _T_14645 = _T_14644 & addrKnown_1; // @[LoadQueue.scala 152:41:@15059.4]
  assign _T_14646 = addrQ_1 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15060.4]
  assign conflict_1_9 = _T_14645 & _T_14646; // @[LoadQueue.scala 152:68:@15061.4]
  assign _T_14648 = entriesToCheck_1_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15063.4]
  assign _T_14649 = _T_14648 & addrKnown_1; // @[LoadQueue.scala 152:41:@15064.4]
  assign _T_14650 = addrQ_1 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15065.4]
  assign conflict_1_10 = _T_14649 & _T_14650; // @[LoadQueue.scala 152:68:@15066.4]
  assign _T_14652 = entriesToCheck_1_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15068.4]
  assign _T_14653 = _T_14652 & addrKnown_1; // @[LoadQueue.scala 152:41:@15069.4]
  assign _T_14654 = addrQ_1 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15070.4]
  assign conflict_1_11 = _T_14653 & _T_14654; // @[LoadQueue.scala 152:68:@15071.4]
  assign _T_14656 = entriesToCheck_1_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15073.4]
  assign _T_14657 = _T_14656 & addrKnown_1; // @[LoadQueue.scala 152:41:@15074.4]
  assign _T_14658 = addrQ_1 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15075.4]
  assign conflict_1_12 = _T_14657 & _T_14658; // @[LoadQueue.scala 152:68:@15076.4]
  assign _T_14660 = entriesToCheck_1_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15078.4]
  assign _T_14661 = _T_14660 & addrKnown_1; // @[LoadQueue.scala 152:41:@15079.4]
  assign _T_14662 = addrQ_1 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15080.4]
  assign conflict_1_13 = _T_14661 & _T_14662; // @[LoadQueue.scala 152:68:@15081.4]
  assign _T_14664 = entriesToCheck_1_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15083.4]
  assign _T_14665 = _T_14664 & addrKnown_1; // @[LoadQueue.scala 152:41:@15084.4]
  assign _T_14666 = addrQ_1 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15085.4]
  assign conflict_1_14 = _T_14665 & _T_14666; // @[LoadQueue.scala 152:68:@15086.4]
  assign _T_14668 = entriesToCheck_1_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15088.4]
  assign _T_14669 = _T_14668 & addrKnown_1; // @[LoadQueue.scala 152:41:@15089.4]
  assign _T_14670 = addrQ_1 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15090.4]
  assign conflict_1_15 = _T_14669 & _T_14670; // @[LoadQueue.scala 152:68:@15091.4]
  assign _T_14672 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15093.4]
  assign _T_14673 = _T_14672 & addrKnown_2; // @[LoadQueue.scala 152:41:@15094.4]
  assign _T_14674 = addrQ_2 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15095.4]
  assign conflict_2_0 = _T_14673 & _T_14674; // @[LoadQueue.scala 152:68:@15096.4]
  assign _T_14676 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15098.4]
  assign _T_14677 = _T_14676 & addrKnown_2; // @[LoadQueue.scala 152:41:@15099.4]
  assign _T_14678 = addrQ_2 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15100.4]
  assign conflict_2_1 = _T_14677 & _T_14678; // @[LoadQueue.scala 152:68:@15101.4]
  assign _T_14680 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15103.4]
  assign _T_14681 = _T_14680 & addrKnown_2; // @[LoadQueue.scala 152:41:@15104.4]
  assign _T_14682 = addrQ_2 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15105.4]
  assign conflict_2_2 = _T_14681 & _T_14682; // @[LoadQueue.scala 152:68:@15106.4]
  assign _T_14684 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15108.4]
  assign _T_14685 = _T_14684 & addrKnown_2; // @[LoadQueue.scala 152:41:@15109.4]
  assign _T_14686 = addrQ_2 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15110.4]
  assign conflict_2_3 = _T_14685 & _T_14686; // @[LoadQueue.scala 152:68:@15111.4]
  assign _T_14688 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15113.4]
  assign _T_14689 = _T_14688 & addrKnown_2; // @[LoadQueue.scala 152:41:@15114.4]
  assign _T_14690 = addrQ_2 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15115.4]
  assign conflict_2_4 = _T_14689 & _T_14690; // @[LoadQueue.scala 152:68:@15116.4]
  assign _T_14692 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15118.4]
  assign _T_14693 = _T_14692 & addrKnown_2; // @[LoadQueue.scala 152:41:@15119.4]
  assign _T_14694 = addrQ_2 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15120.4]
  assign conflict_2_5 = _T_14693 & _T_14694; // @[LoadQueue.scala 152:68:@15121.4]
  assign _T_14696 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15123.4]
  assign _T_14697 = _T_14696 & addrKnown_2; // @[LoadQueue.scala 152:41:@15124.4]
  assign _T_14698 = addrQ_2 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15125.4]
  assign conflict_2_6 = _T_14697 & _T_14698; // @[LoadQueue.scala 152:68:@15126.4]
  assign _T_14700 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15128.4]
  assign _T_14701 = _T_14700 & addrKnown_2; // @[LoadQueue.scala 152:41:@15129.4]
  assign _T_14702 = addrQ_2 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15130.4]
  assign conflict_2_7 = _T_14701 & _T_14702; // @[LoadQueue.scala 152:68:@15131.4]
  assign _T_14704 = entriesToCheck_2_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15133.4]
  assign _T_14705 = _T_14704 & addrKnown_2; // @[LoadQueue.scala 152:41:@15134.4]
  assign _T_14706 = addrQ_2 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15135.4]
  assign conflict_2_8 = _T_14705 & _T_14706; // @[LoadQueue.scala 152:68:@15136.4]
  assign _T_14708 = entriesToCheck_2_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15138.4]
  assign _T_14709 = _T_14708 & addrKnown_2; // @[LoadQueue.scala 152:41:@15139.4]
  assign _T_14710 = addrQ_2 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15140.4]
  assign conflict_2_9 = _T_14709 & _T_14710; // @[LoadQueue.scala 152:68:@15141.4]
  assign _T_14712 = entriesToCheck_2_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15143.4]
  assign _T_14713 = _T_14712 & addrKnown_2; // @[LoadQueue.scala 152:41:@15144.4]
  assign _T_14714 = addrQ_2 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15145.4]
  assign conflict_2_10 = _T_14713 & _T_14714; // @[LoadQueue.scala 152:68:@15146.4]
  assign _T_14716 = entriesToCheck_2_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15148.4]
  assign _T_14717 = _T_14716 & addrKnown_2; // @[LoadQueue.scala 152:41:@15149.4]
  assign _T_14718 = addrQ_2 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15150.4]
  assign conflict_2_11 = _T_14717 & _T_14718; // @[LoadQueue.scala 152:68:@15151.4]
  assign _T_14720 = entriesToCheck_2_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15153.4]
  assign _T_14721 = _T_14720 & addrKnown_2; // @[LoadQueue.scala 152:41:@15154.4]
  assign _T_14722 = addrQ_2 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15155.4]
  assign conflict_2_12 = _T_14721 & _T_14722; // @[LoadQueue.scala 152:68:@15156.4]
  assign _T_14724 = entriesToCheck_2_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15158.4]
  assign _T_14725 = _T_14724 & addrKnown_2; // @[LoadQueue.scala 152:41:@15159.4]
  assign _T_14726 = addrQ_2 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15160.4]
  assign conflict_2_13 = _T_14725 & _T_14726; // @[LoadQueue.scala 152:68:@15161.4]
  assign _T_14728 = entriesToCheck_2_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15163.4]
  assign _T_14729 = _T_14728 & addrKnown_2; // @[LoadQueue.scala 152:41:@15164.4]
  assign _T_14730 = addrQ_2 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15165.4]
  assign conflict_2_14 = _T_14729 & _T_14730; // @[LoadQueue.scala 152:68:@15166.4]
  assign _T_14732 = entriesToCheck_2_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15168.4]
  assign _T_14733 = _T_14732 & addrKnown_2; // @[LoadQueue.scala 152:41:@15169.4]
  assign _T_14734 = addrQ_2 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15170.4]
  assign conflict_2_15 = _T_14733 & _T_14734; // @[LoadQueue.scala 152:68:@15171.4]
  assign _T_14736 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15173.4]
  assign _T_14737 = _T_14736 & addrKnown_3; // @[LoadQueue.scala 152:41:@15174.4]
  assign _T_14738 = addrQ_3 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15175.4]
  assign conflict_3_0 = _T_14737 & _T_14738; // @[LoadQueue.scala 152:68:@15176.4]
  assign _T_14740 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15178.4]
  assign _T_14741 = _T_14740 & addrKnown_3; // @[LoadQueue.scala 152:41:@15179.4]
  assign _T_14742 = addrQ_3 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15180.4]
  assign conflict_3_1 = _T_14741 & _T_14742; // @[LoadQueue.scala 152:68:@15181.4]
  assign _T_14744 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15183.4]
  assign _T_14745 = _T_14744 & addrKnown_3; // @[LoadQueue.scala 152:41:@15184.4]
  assign _T_14746 = addrQ_3 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15185.4]
  assign conflict_3_2 = _T_14745 & _T_14746; // @[LoadQueue.scala 152:68:@15186.4]
  assign _T_14748 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15188.4]
  assign _T_14749 = _T_14748 & addrKnown_3; // @[LoadQueue.scala 152:41:@15189.4]
  assign _T_14750 = addrQ_3 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15190.4]
  assign conflict_3_3 = _T_14749 & _T_14750; // @[LoadQueue.scala 152:68:@15191.4]
  assign _T_14752 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15193.4]
  assign _T_14753 = _T_14752 & addrKnown_3; // @[LoadQueue.scala 152:41:@15194.4]
  assign _T_14754 = addrQ_3 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15195.4]
  assign conflict_3_4 = _T_14753 & _T_14754; // @[LoadQueue.scala 152:68:@15196.4]
  assign _T_14756 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15198.4]
  assign _T_14757 = _T_14756 & addrKnown_3; // @[LoadQueue.scala 152:41:@15199.4]
  assign _T_14758 = addrQ_3 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15200.4]
  assign conflict_3_5 = _T_14757 & _T_14758; // @[LoadQueue.scala 152:68:@15201.4]
  assign _T_14760 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15203.4]
  assign _T_14761 = _T_14760 & addrKnown_3; // @[LoadQueue.scala 152:41:@15204.4]
  assign _T_14762 = addrQ_3 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15205.4]
  assign conflict_3_6 = _T_14761 & _T_14762; // @[LoadQueue.scala 152:68:@15206.4]
  assign _T_14764 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15208.4]
  assign _T_14765 = _T_14764 & addrKnown_3; // @[LoadQueue.scala 152:41:@15209.4]
  assign _T_14766 = addrQ_3 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15210.4]
  assign conflict_3_7 = _T_14765 & _T_14766; // @[LoadQueue.scala 152:68:@15211.4]
  assign _T_14768 = entriesToCheck_3_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15213.4]
  assign _T_14769 = _T_14768 & addrKnown_3; // @[LoadQueue.scala 152:41:@15214.4]
  assign _T_14770 = addrQ_3 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15215.4]
  assign conflict_3_8 = _T_14769 & _T_14770; // @[LoadQueue.scala 152:68:@15216.4]
  assign _T_14772 = entriesToCheck_3_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15218.4]
  assign _T_14773 = _T_14772 & addrKnown_3; // @[LoadQueue.scala 152:41:@15219.4]
  assign _T_14774 = addrQ_3 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15220.4]
  assign conflict_3_9 = _T_14773 & _T_14774; // @[LoadQueue.scala 152:68:@15221.4]
  assign _T_14776 = entriesToCheck_3_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15223.4]
  assign _T_14777 = _T_14776 & addrKnown_3; // @[LoadQueue.scala 152:41:@15224.4]
  assign _T_14778 = addrQ_3 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15225.4]
  assign conflict_3_10 = _T_14777 & _T_14778; // @[LoadQueue.scala 152:68:@15226.4]
  assign _T_14780 = entriesToCheck_3_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15228.4]
  assign _T_14781 = _T_14780 & addrKnown_3; // @[LoadQueue.scala 152:41:@15229.4]
  assign _T_14782 = addrQ_3 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15230.4]
  assign conflict_3_11 = _T_14781 & _T_14782; // @[LoadQueue.scala 152:68:@15231.4]
  assign _T_14784 = entriesToCheck_3_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15233.4]
  assign _T_14785 = _T_14784 & addrKnown_3; // @[LoadQueue.scala 152:41:@15234.4]
  assign _T_14786 = addrQ_3 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15235.4]
  assign conflict_3_12 = _T_14785 & _T_14786; // @[LoadQueue.scala 152:68:@15236.4]
  assign _T_14788 = entriesToCheck_3_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15238.4]
  assign _T_14789 = _T_14788 & addrKnown_3; // @[LoadQueue.scala 152:41:@15239.4]
  assign _T_14790 = addrQ_3 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15240.4]
  assign conflict_3_13 = _T_14789 & _T_14790; // @[LoadQueue.scala 152:68:@15241.4]
  assign _T_14792 = entriesToCheck_3_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15243.4]
  assign _T_14793 = _T_14792 & addrKnown_3; // @[LoadQueue.scala 152:41:@15244.4]
  assign _T_14794 = addrQ_3 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15245.4]
  assign conflict_3_14 = _T_14793 & _T_14794; // @[LoadQueue.scala 152:68:@15246.4]
  assign _T_14796 = entriesToCheck_3_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15248.4]
  assign _T_14797 = _T_14796 & addrKnown_3; // @[LoadQueue.scala 152:41:@15249.4]
  assign _T_14798 = addrQ_3 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15250.4]
  assign conflict_3_15 = _T_14797 & _T_14798; // @[LoadQueue.scala 152:68:@15251.4]
  assign _T_14800 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15253.4]
  assign _T_14801 = _T_14800 & addrKnown_4; // @[LoadQueue.scala 152:41:@15254.4]
  assign _T_14802 = addrQ_4 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15255.4]
  assign conflict_4_0 = _T_14801 & _T_14802; // @[LoadQueue.scala 152:68:@15256.4]
  assign _T_14804 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15258.4]
  assign _T_14805 = _T_14804 & addrKnown_4; // @[LoadQueue.scala 152:41:@15259.4]
  assign _T_14806 = addrQ_4 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15260.4]
  assign conflict_4_1 = _T_14805 & _T_14806; // @[LoadQueue.scala 152:68:@15261.4]
  assign _T_14808 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15263.4]
  assign _T_14809 = _T_14808 & addrKnown_4; // @[LoadQueue.scala 152:41:@15264.4]
  assign _T_14810 = addrQ_4 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15265.4]
  assign conflict_4_2 = _T_14809 & _T_14810; // @[LoadQueue.scala 152:68:@15266.4]
  assign _T_14812 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15268.4]
  assign _T_14813 = _T_14812 & addrKnown_4; // @[LoadQueue.scala 152:41:@15269.4]
  assign _T_14814 = addrQ_4 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15270.4]
  assign conflict_4_3 = _T_14813 & _T_14814; // @[LoadQueue.scala 152:68:@15271.4]
  assign _T_14816 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15273.4]
  assign _T_14817 = _T_14816 & addrKnown_4; // @[LoadQueue.scala 152:41:@15274.4]
  assign _T_14818 = addrQ_4 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15275.4]
  assign conflict_4_4 = _T_14817 & _T_14818; // @[LoadQueue.scala 152:68:@15276.4]
  assign _T_14820 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15278.4]
  assign _T_14821 = _T_14820 & addrKnown_4; // @[LoadQueue.scala 152:41:@15279.4]
  assign _T_14822 = addrQ_4 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15280.4]
  assign conflict_4_5 = _T_14821 & _T_14822; // @[LoadQueue.scala 152:68:@15281.4]
  assign _T_14824 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15283.4]
  assign _T_14825 = _T_14824 & addrKnown_4; // @[LoadQueue.scala 152:41:@15284.4]
  assign _T_14826 = addrQ_4 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15285.4]
  assign conflict_4_6 = _T_14825 & _T_14826; // @[LoadQueue.scala 152:68:@15286.4]
  assign _T_14828 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15288.4]
  assign _T_14829 = _T_14828 & addrKnown_4; // @[LoadQueue.scala 152:41:@15289.4]
  assign _T_14830 = addrQ_4 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15290.4]
  assign conflict_4_7 = _T_14829 & _T_14830; // @[LoadQueue.scala 152:68:@15291.4]
  assign _T_14832 = entriesToCheck_4_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15293.4]
  assign _T_14833 = _T_14832 & addrKnown_4; // @[LoadQueue.scala 152:41:@15294.4]
  assign _T_14834 = addrQ_4 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15295.4]
  assign conflict_4_8 = _T_14833 & _T_14834; // @[LoadQueue.scala 152:68:@15296.4]
  assign _T_14836 = entriesToCheck_4_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15298.4]
  assign _T_14837 = _T_14836 & addrKnown_4; // @[LoadQueue.scala 152:41:@15299.4]
  assign _T_14838 = addrQ_4 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15300.4]
  assign conflict_4_9 = _T_14837 & _T_14838; // @[LoadQueue.scala 152:68:@15301.4]
  assign _T_14840 = entriesToCheck_4_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15303.4]
  assign _T_14841 = _T_14840 & addrKnown_4; // @[LoadQueue.scala 152:41:@15304.4]
  assign _T_14842 = addrQ_4 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15305.4]
  assign conflict_4_10 = _T_14841 & _T_14842; // @[LoadQueue.scala 152:68:@15306.4]
  assign _T_14844 = entriesToCheck_4_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15308.4]
  assign _T_14845 = _T_14844 & addrKnown_4; // @[LoadQueue.scala 152:41:@15309.4]
  assign _T_14846 = addrQ_4 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15310.4]
  assign conflict_4_11 = _T_14845 & _T_14846; // @[LoadQueue.scala 152:68:@15311.4]
  assign _T_14848 = entriesToCheck_4_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15313.4]
  assign _T_14849 = _T_14848 & addrKnown_4; // @[LoadQueue.scala 152:41:@15314.4]
  assign _T_14850 = addrQ_4 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15315.4]
  assign conflict_4_12 = _T_14849 & _T_14850; // @[LoadQueue.scala 152:68:@15316.4]
  assign _T_14852 = entriesToCheck_4_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15318.4]
  assign _T_14853 = _T_14852 & addrKnown_4; // @[LoadQueue.scala 152:41:@15319.4]
  assign _T_14854 = addrQ_4 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15320.4]
  assign conflict_4_13 = _T_14853 & _T_14854; // @[LoadQueue.scala 152:68:@15321.4]
  assign _T_14856 = entriesToCheck_4_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15323.4]
  assign _T_14857 = _T_14856 & addrKnown_4; // @[LoadQueue.scala 152:41:@15324.4]
  assign _T_14858 = addrQ_4 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15325.4]
  assign conflict_4_14 = _T_14857 & _T_14858; // @[LoadQueue.scala 152:68:@15326.4]
  assign _T_14860 = entriesToCheck_4_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15328.4]
  assign _T_14861 = _T_14860 & addrKnown_4; // @[LoadQueue.scala 152:41:@15329.4]
  assign _T_14862 = addrQ_4 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15330.4]
  assign conflict_4_15 = _T_14861 & _T_14862; // @[LoadQueue.scala 152:68:@15331.4]
  assign _T_14864 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15333.4]
  assign _T_14865 = _T_14864 & addrKnown_5; // @[LoadQueue.scala 152:41:@15334.4]
  assign _T_14866 = addrQ_5 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15335.4]
  assign conflict_5_0 = _T_14865 & _T_14866; // @[LoadQueue.scala 152:68:@15336.4]
  assign _T_14868 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15338.4]
  assign _T_14869 = _T_14868 & addrKnown_5; // @[LoadQueue.scala 152:41:@15339.4]
  assign _T_14870 = addrQ_5 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15340.4]
  assign conflict_5_1 = _T_14869 & _T_14870; // @[LoadQueue.scala 152:68:@15341.4]
  assign _T_14872 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15343.4]
  assign _T_14873 = _T_14872 & addrKnown_5; // @[LoadQueue.scala 152:41:@15344.4]
  assign _T_14874 = addrQ_5 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15345.4]
  assign conflict_5_2 = _T_14873 & _T_14874; // @[LoadQueue.scala 152:68:@15346.4]
  assign _T_14876 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15348.4]
  assign _T_14877 = _T_14876 & addrKnown_5; // @[LoadQueue.scala 152:41:@15349.4]
  assign _T_14878 = addrQ_5 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15350.4]
  assign conflict_5_3 = _T_14877 & _T_14878; // @[LoadQueue.scala 152:68:@15351.4]
  assign _T_14880 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15353.4]
  assign _T_14881 = _T_14880 & addrKnown_5; // @[LoadQueue.scala 152:41:@15354.4]
  assign _T_14882 = addrQ_5 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15355.4]
  assign conflict_5_4 = _T_14881 & _T_14882; // @[LoadQueue.scala 152:68:@15356.4]
  assign _T_14884 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15358.4]
  assign _T_14885 = _T_14884 & addrKnown_5; // @[LoadQueue.scala 152:41:@15359.4]
  assign _T_14886 = addrQ_5 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15360.4]
  assign conflict_5_5 = _T_14885 & _T_14886; // @[LoadQueue.scala 152:68:@15361.4]
  assign _T_14888 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15363.4]
  assign _T_14889 = _T_14888 & addrKnown_5; // @[LoadQueue.scala 152:41:@15364.4]
  assign _T_14890 = addrQ_5 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15365.4]
  assign conflict_5_6 = _T_14889 & _T_14890; // @[LoadQueue.scala 152:68:@15366.4]
  assign _T_14892 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15368.4]
  assign _T_14893 = _T_14892 & addrKnown_5; // @[LoadQueue.scala 152:41:@15369.4]
  assign _T_14894 = addrQ_5 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15370.4]
  assign conflict_5_7 = _T_14893 & _T_14894; // @[LoadQueue.scala 152:68:@15371.4]
  assign _T_14896 = entriesToCheck_5_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15373.4]
  assign _T_14897 = _T_14896 & addrKnown_5; // @[LoadQueue.scala 152:41:@15374.4]
  assign _T_14898 = addrQ_5 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15375.4]
  assign conflict_5_8 = _T_14897 & _T_14898; // @[LoadQueue.scala 152:68:@15376.4]
  assign _T_14900 = entriesToCheck_5_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15378.4]
  assign _T_14901 = _T_14900 & addrKnown_5; // @[LoadQueue.scala 152:41:@15379.4]
  assign _T_14902 = addrQ_5 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15380.4]
  assign conflict_5_9 = _T_14901 & _T_14902; // @[LoadQueue.scala 152:68:@15381.4]
  assign _T_14904 = entriesToCheck_5_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15383.4]
  assign _T_14905 = _T_14904 & addrKnown_5; // @[LoadQueue.scala 152:41:@15384.4]
  assign _T_14906 = addrQ_5 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15385.4]
  assign conflict_5_10 = _T_14905 & _T_14906; // @[LoadQueue.scala 152:68:@15386.4]
  assign _T_14908 = entriesToCheck_5_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15388.4]
  assign _T_14909 = _T_14908 & addrKnown_5; // @[LoadQueue.scala 152:41:@15389.4]
  assign _T_14910 = addrQ_5 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15390.4]
  assign conflict_5_11 = _T_14909 & _T_14910; // @[LoadQueue.scala 152:68:@15391.4]
  assign _T_14912 = entriesToCheck_5_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15393.4]
  assign _T_14913 = _T_14912 & addrKnown_5; // @[LoadQueue.scala 152:41:@15394.4]
  assign _T_14914 = addrQ_5 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15395.4]
  assign conflict_5_12 = _T_14913 & _T_14914; // @[LoadQueue.scala 152:68:@15396.4]
  assign _T_14916 = entriesToCheck_5_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15398.4]
  assign _T_14917 = _T_14916 & addrKnown_5; // @[LoadQueue.scala 152:41:@15399.4]
  assign _T_14918 = addrQ_5 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15400.4]
  assign conflict_5_13 = _T_14917 & _T_14918; // @[LoadQueue.scala 152:68:@15401.4]
  assign _T_14920 = entriesToCheck_5_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15403.4]
  assign _T_14921 = _T_14920 & addrKnown_5; // @[LoadQueue.scala 152:41:@15404.4]
  assign _T_14922 = addrQ_5 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15405.4]
  assign conflict_5_14 = _T_14921 & _T_14922; // @[LoadQueue.scala 152:68:@15406.4]
  assign _T_14924 = entriesToCheck_5_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15408.4]
  assign _T_14925 = _T_14924 & addrKnown_5; // @[LoadQueue.scala 152:41:@15409.4]
  assign _T_14926 = addrQ_5 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15410.4]
  assign conflict_5_15 = _T_14925 & _T_14926; // @[LoadQueue.scala 152:68:@15411.4]
  assign _T_14928 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15413.4]
  assign _T_14929 = _T_14928 & addrKnown_6; // @[LoadQueue.scala 152:41:@15414.4]
  assign _T_14930 = addrQ_6 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15415.4]
  assign conflict_6_0 = _T_14929 & _T_14930; // @[LoadQueue.scala 152:68:@15416.4]
  assign _T_14932 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15418.4]
  assign _T_14933 = _T_14932 & addrKnown_6; // @[LoadQueue.scala 152:41:@15419.4]
  assign _T_14934 = addrQ_6 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15420.4]
  assign conflict_6_1 = _T_14933 & _T_14934; // @[LoadQueue.scala 152:68:@15421.4]
  assign _T_14936 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15423.4]
  assign _T_14937 = _T_14936 & addrKnown_6; // @[LoadQueue.scala 152:41:@15424.4]
  assign _T_14938 = addrQ_6 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15425.4]
  assign conflict_6_2 = _T_14937 & _T_14938; // @[LoadQueue.scala 152:68:@15426.4]
  assign _T_14940 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15428.4]
  assign _T_14941 = _T_14940 & addrKnown_6; // @[LoadQueue.scala 152:41:@15429.4]
  assign _T_14942 = addrQ_6 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15430.4]
  assign conflict_6_3 = _T_14941 & _T_14942; // @[LoadQueue.scala 152:68:@15431.4]
  assign _T_14944 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15433.4]
  assign _T_14945 = _T_14944 & addrKnown_6; // @[LoadQueue.scala 152:41:@15434.4]
  assign _T_14946 = addrQ_6 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15435.4]
  assign conflict_6_4 = _T_14945 & _T_14946; // @[LoadQueue.scala 152:68:@15436.4]
  assign _T_14948 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15438.4]
  assign _T_14949 = _T_14948 & addrKnown_6; // @[LoadQueue.scala 152:41:@15439.4]
  assign _T_14950 = addrQ_6 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15440.4]
  assign conflict_6_5 = _T_14949 & _T_14950; // @[LoadQueue.scala 152:68:@15441.4]
  assign _T_14952 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15443.4]
  assign _T_14953 = _T_14952 & addrKnown_6; // @[LoadQueue.scala 152:41:@15444.4]
  assign _T_14954 = addrQ_6 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15445.4]
  assign conflict_6_6 = _T_14953 & _T_14954; // @[LoadQueue.scala 152:68:@15446.4]
  assign _T_14956 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15448.4]
  assign _T_14957 = _T_14956 & addrKnown_6; // @[LoadQueue.scala 152:41:@15449.4]
  assign _T_14958 = addrQ_6 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15450.4]
  assign conflict_6_7 = _T_14957 & _T_14958; // @[LoadQueue.scala 152:68:@15451.4]
  assign _T_14960 = entriesToCheck_6_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15453.4]
  assign _T_14961 = _T_14960 & addrKnown_6; // @[LoadQueue.scala 152:41:@15454.4]
  assign _T_14962 = addrQ_6 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15455.4]
  assign conflict_6_8 = _T_14961 & _T_14962; // @[LoadQueue.scala 152:68:@15456.4]
  assign _T_14964 = entriesToCheck_6_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15458.4]
  assign _T_14965 = _T_14964 & addrKnown_6; // @[LoadQueue.scala 152:41:@15459.4]
  assign _T_14966 = addrQ_6 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15460.4]
  assign conflict_6_9 = _T_14965 & _T_14966; // @[LoadQueue.scala 152:68:@15461.4]
  assign _T_14968 = entriesToCheck_6_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15463.4]
  assign _T_14969 = _T_14968 & addrKnown_6; // @[LoadQueue.scala 152:41:@15464.4]
  assign _T_14970 = addrQ_6 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15465.4]
  assign conflict_6_10 = _T_14969 & _T_14970; // @[LoadQueue.scala 152:68:@15466.4]
  assign _T_14972 = entriesToCheck_6_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15468.4]
  assign _T_14973 = _T_14972 & addrKnown_6; // @[LoadQueue.scala 152:41:@15469.4]
  assign _T_14974 = addrQ_6 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15470.4]
  assign conflict_6_11 = _T_14973 & _T_14974; // @[LoadQueue.scala 152:68:@15471.4]
  assign _T_14976 = entriesToCheck_6_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15473.4]
  assign _T_14977 = _T_14976 & addrKnown_6; // @[LoadQueue.scala 152:41:@15474.4]
  assign _T_14978 = addrQ_6 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15475.4]
  assign conflict_6_12 = _T_14977 & _T_14978; // @[LoadQueue.scala 152:68:@15476.4]
  assign _T_14980 = entriesToCheck_6_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15478.4]
  assign _T_14981 = _T_14980 & addrKnown_6; // @[LoadQueue.scala 152:41:@15479.4]
  assign _T_14982 = addrQ_6 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15480.4]
  assign conflict_6_13 = _T_14981 & _T_14982; // @[LoadQueue.scala 152:68:@15481.4]
  assign _T_14984 = entriesToCheck_6_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15483.4]
  assign _T_14985 = _T_14984 & addrKnown_6; // @[LoadQueue.scala 152:41:@15484.4]
  assign _T_14986 = addrQ_6 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15485.4]
  assign conflict_6_14 = _T_14985 & _T_14986; // @[LoadQueue.scala 152:68:@15486.4]
  assign _T_14988 = entriesToCheck_6_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15488.4]
  assign _T_14989 = _T_14988 & addrKnown_6; // @[LoadQueue.scala 152:41:@15489.4]
  assign _T_14990 = addrQ_6 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15490.4]
  assign conflict_6_15 = _T_14989 & _T_14990; // @[LoadQueue.scala 152:68:@15491.4]
  assign _T_14992 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15493.4]
  assign _T_14993 = _T_14992 & addrKnown_7; // @[LoadQueue.scala 152:41:@15494.4]
  assign _T_14994 = addrQ_7 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15495.4]
  assign conflict_7_0 = _T_14993 & _T_14994; // @[LoadQueue.scala 152:68:@15496.4]
  assign _T_14996 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15498.4]
  assign _T_14997 = _T_14996 & addrKnown_7; // @[LoadQueue.scala 152:41:@15499.4]
  assign _T_14998 = addrQ_7 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15500.4]
  assign conflict_7_1 = _T_14997 & _T_14998; // @[LoadQueue.scala 152:68:@15501.4]
  assign _T_15000 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15503.4]
  assign _T_15001 = _T_15000 & addrKnown_7; // @[LoadQueue.scala 152:41:@15504.4]
  assign _T_15002 = addrQ_7 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15505.4]
  assign conflict_7_2 = _T_15001 & _T_15002; // @[LoadQueue.scala 152:68:@15506.4]
  assign _T_15004 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15508.4]
  assign _T_15005 = _T_15004 & addrKnown_7; // @[LoadQueue.scala 152:41:@15509.4]
  assign _T_15006 = addrQ_7 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15510.4]
  assign conflict_7_3 = _T_15005 & _T_15006; // @[LoadQueue.scala 152:68:@15511.4]
  assign _T_15008 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15513.4]
  assign _T_15009 = _T_15008 & addrKnown_7; // @[LoadQueue.scala 152:41:@15514.4]
  assign _T_15010 = addrQ_7 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15515.4]
  assign conflict_7_4 = _T_15009 & _T_15010; // @[LoadQueue.scala 152:68:@15516.4]
  assign _T_15012 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15518.4]
  assign _T_15013 = _T_15012 & addrKnown_7; // @[LoadQueue.scala 152:41:@15519.4]
  assign _T_15014 = addrQ_7 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15520.4]
  assign conflict_7_5 = _T_15013 & _T_15014; // @[LoadQueue.scala 152:68:@15521.4]
  assign _T_15016 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15523.4]
  assign _T_15017 = _T_15016 & addrKnown_7; // @[LoadQueue.scala 152:41:@15524.4]
  assign _T_15018 = addrQ_7 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15525.4]
  assign conflict_7_6 = _T_15017 & _T_15018; // @[LoadQueue.scala 152:68:@15526.4]
  assign _T_15020 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15528.4]
  assign _T_15021 = _T_15020 & addrKnown_7; // @[LoadQueue.scala 152:41:@15529.4]
  assign _T_15022 = addrQ_7 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15530.4]
  assign conflict_7_7 = _T_15021 & _T_15022; // @[LoadQueue.scala 152:68:@15531.4]
  assign _T_15024 = entriesToCheck_7_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15533.4]
  assign _T_15025 = _T_15024 & addrKnown_7; // @[LoadQueue.scala 152:41:@15534.4]
  assign _T_15026 = addrQ_7 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15535.4]
  assign conflict_7_8 = _T_15025 & _T_15026; // @[LoadQueue.scala 152:68:@15536.4]
  assign _T_15028 = entriesToCheck_7_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15538.4]
  assign _T_15029 = _T_15028 & addrKnown_7; // @[LoadQueue.scala 152:41:@15539.4]
  assign _T_15030 = addrQ_7 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15540.4]
  assign conflict_7_9 = _T_15029 & _T_15030; // @[LoadQueue.scala 152:68:@15541.4]
  assign _T_15032 = entriesToCheck_7_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15543.4]
  assign _T_15033 = _T_15032 & addrKnown_7; // @[LoadQueue.scala 152:41:@15544.4]
  assign _T_15034 = addrQ_7 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15545.4]
  assign conflict_7_10 = _T_15033 & _T_15034; // @[LoadQueue.scala 152:68:@15546.4]
  assign _T_15036 = entriesToCheck_7_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15548.4]
  assign _T_15037 = _T_15036 & addrKnown_7; // @[LoadQueue.scala 152:41:@15549.4]
  assign _T_15038 = addrQ_7 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15550.4]
  assign conflict_7_11 = _T_15037 & _T_15038; // @[LoadQueue.scala 152:68:@15551.4]
  assign _T_15040 = entriesToCheck_7_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15553.4]
  assign _T_15041 = _T_15040 & addrKnown_7; // @[LoadQueue.scala 152:41:@15554.4]
  assign _T_15042 = addrQ_7 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15555.4]
  assign conflict_7_12 = _T_15041 & _T_15042; // @[LoadQueue.scala 152:68:@15556.4]
  assign _T_15044 = entriesToCheck_7_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15558.4]
  assign _T_15045 = _T_15044 & addrKnown_7; // @[LoadQueue.scala 152:41:@15559.4]
  assign _T_15046 = addrQ_7 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15560.4]
  assign conflict_7_13 = _T_15045 & _T_15046; // @[LoadQueue.scala 152:68:@15561.4]
  assign _T_15048 = entriesToCheck_7_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15563.4]
  assign _T_15049 = _T_15048 & addrKnown_7; // @[LoadQueue.scala 152:41:@15564.4]
  assign _T_15050 = addrQ_7 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15565.4]
  assign conflict_7_14 = _T_15049 & _T_15050; // @[LoadQueue.scala 152:68:@15566.4]
  assign _T_15052 = entriesToCheck_7_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15568.4]
  assign _T_15053 = _T_15052 & addrKnown_7; // @[LoadQueue.scala 152:41:@15569.4]
  assign _T_15054 = addrQ_7 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15570.4]
  assign conflict_7_15 = _T_15053 & _T_15054; // @[LoadQueue.scala 152:68:@15571.4]
  assign _T_15056 = entriesToCheck_8_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15573.4]
  assign _T_15057 = _T_15056 & addrKnown_8; // @[LoadQueue.scala 152:41:@15574.4]
  assign _T_15058 = addrQ_8 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15575.4]
  assign conflict_8_0 = _T_15057 & _T_15058; // @[LoadQueue.scala 152:68:@15576.4]
  assign _T_15060 = entriesToCheck_8_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15578.4]
  assign _T_15061 = _T_15060 & addrKnown_8; // @[LoadQueue.scala 152:41:@15579.4]
  assign _T_15062 = addrQ_8 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15580.4]
  assign conflict_8_1 = _T_15061 & _T_15062; // @[LoadQueue.scala 152:68:@15581.4]
  assign _T_15064 = entriesToCheck_8_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15583.4]
  assign _T_15065 = _T_15064 & addrKnown_8; // @[LoadQueue.scala 152:41:@15584.4]
  assign _T_15066 = addrQ_8 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15585.4]
  assign conflict_8_2 = _T_15065 & _T_15066; // @[LoadQueue.scala 152:68:@15586.4]
  assign _T_15068 = entriesToCheck_8_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15588.4]
  assign _T_15069 = _T_15068 & addrKnown_8; // @[LoadQueue.scala 152:41:@15589.4]
  assign _T_15070 = addrQ_8 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15590.4]
  assign conflict_8_3 = _T_15069 & _T_15070; // @[LoadQueue.scala 152:68:@15591.4]
  assign _T_15072 = entriesToCheck_8_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15593.4]
  assign _T_15073 = _T_15072 & addrKnown_8; // @[LoadQueue.scala 152:41:@15594.4]
  assign _T_15074 = addrQ_8 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15595.4]
  assign conflict_8_4 = _T_15073 & _T_15074; // @[LoadQueue.scala 152:68:@15596.4]
  assign _T_15076 = entriesToCheck_8_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15598.4]
  assign _T_15077 = _T_15076 & addrKnown_8; // @[LoadQueue.scala 152:41:@15599.4]
  assign _T_15078 = addrQ_8 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15600.4]
  assign conflict_8_5 = _T_15077 & _T_15078; // @[LoadQueue.scala 152:68:@15601.4]
  assign _T_15080 = entriesToCheck_8_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15603.4]
  assign _T_15081 = _T_15080 & addrKnown_8; // @[LoadQueue.scala 152:41:@15604.4]
  assign _T_15082 = addrQ_8 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15605.4]
  assign conflict_8_6 = _T_15081 & _T_15082; // @[LoadQueue.scala 152:68:@15606.4]
  assign _T_15084 = entriesToCheck_8_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15608.4]
  assign _T_15085 = _T_15084 & addrKnown_8; // @[LoadQueue.scala 152:41:@15609.4]
  assign _T_15086 = addrQ_8 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15610.4]
  assign conflict_8_7 = _T_15085 & _T_15086; // @[LoadQueue.scala 152:68:@15611.4]
  assign _T_15088 = entriesToCheck_8_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15613.4]
  assign _T_15089 = _T_15088 & addrKnown_8; // @[LoadQueue.scala 152:41:@15614.4]
  assign _T_15090 = addrQ_8 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15615.4]
  assign conflict_8_8 = _T_15089 & _T_15090; // @[LoadQueue.scala 152:68:@15616.4]
  assign _T_15092 = entriesToCheck_8_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15618.4]
  assign _T_15093 = _T_15092 & addrKnown_8; // @[LoadQueue.scala 152:41:@15619.4]
  assign _T_15094 = addrQ_8 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15620.4]
  assign conflict_8_9 = _T_15093 & _T_15094; // @[LoadQueue.scala 152:68:@15621.4]
  assign _T_15096 = entriesToCheck_8_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15623.4]
  assign _T_15097 = _T_15096 & addrKnown_8; // @[LoadQueue.scala 152:41:@15624.4]
  assign _T_15098 = addrQ_8 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15625.4]
  assign conflict_8_10 = _T_15097 & _T_15098; // @[LoadQueue.scala 152:68:@15626.4]
  assign _T_15100 = entriesToCheck_8_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15628.4]
  assign _T_15101 = _T_15100 & addrKnown_8; // @[LoadQueue.scala 152:41:@15629.4]
  assign _T_15102 = addrQ_8 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15630.4]
  assign conflict_8_11 = _T_15101 & _T_15102; // @[LoadQueue.scala 152:68:@15631.4]
  assign _T_15104 = entriesToCheck_8_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15633.4]
  assign _T_15105 = _T_15104 & addrKnown_8; // @[LoadQueue.scala 152:41:@15634.4]
  assign _T_15106 = addrQ_8 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15635.4]
  assign conflict_8_12 = _T_15105 & _T_15106; // @[LoadQueue.scala 152:68:@15636.4]
  assign _T_15108 = entriesToCheck_8_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15638.4]
  assign _T_15109 = _T_15108 & addrKnown_8; // @[LoadQueue.scala 152:41:@15639.4]
  assign _T_15110 = addrQ_8 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15640.4]
  assign conflict_8_13 = _T_15109 & _T_15110; // @[LoadQueue.scala 152:68:@15641.4]
  assign _T_15112 = entriesToCheck_8_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15643.4]
  assign _T_15113 = _T_15112 & addrKnown_8; // @[LoadQueue.scala 152:41:@15644.4]
  assign _T_15114 = addrQ_8 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15645.4]
  assign conflict_8_14 = _T_15113 & _T_15114; // @[LoadQueue.scala 152:68:@15646.4]
  assign _T_15116 = entriesToCheck_8_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15648.4]
  assign _T_15117 = _T_15116 & addrKnown_8; // @[LoadQueue.scala 152:41:@15649.4]
  assign _T_15118 = addrQ_8 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15650.4]
  assign conflict_8_15 = _T_15117 & _T_15118; // @[LoadQueue.scala 152:68:@15651.4]
  assign _T_15120 = entriesToCheck_9_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15653.4]
  assign _T_15121 = _T_15120 & addrKnown_9; // @[LoadQueue.scala 152:41:@15654.4]
  assign _T_15122 = addrQ_9 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15655.4]
  assign conflict_9_0 = _T_15121 & _T_15122; // @[LoadQueue.scala 152:68:@15656.4]
  assign _T_15124 = entriesToCheck_9_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15658.4]
  assign _T_15125 = _T_15124 & addrKnown_9; // @[LoadQueue.scala 152:41:@15659.4]
  assign _T_15126 = addrQ_9 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15660.4]
  assign conflict_9_1 = _T_15125 & _T_15126; // @[LoadQueue.scala 152:68:@15661.4]
  assign _T_15128 = entriesToCheck_9_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15663.4]
  assign _T_15129 = _T_15128 & addrKnown_9; // @[LoadQueue.scala 152:41:@15664.4]
  assign _T_15130 = addrQ_9 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15665.4]
  assign conflict_9_2 = _T_15129 & _T_15130; // @[LoadQueue.scala 152:68:@15666.4]
  assign _T_15132 = entriesToCheck_9_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15668.4]
  assign _T_15133 = _T_15132 & addrKnown_9; // @[LoadQueue.scala 152:41:@15669.4]
  assign _T_15134 = addrQ_9 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15670.4]
  assign conflict_9_3 = _T_15133 & _T_15134; // @[LoadQueue.scala 152:68:@15671.4]
  assign _T_15136 = entriesToCheck_9_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15673.4]
  assign _T_15137 = _T_15136 & addrKnown_9; // @[LoadQueue.scala 152:41:@15674.4]
  assign _T_15138 = addrQ_9 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15675.4]
  assign conflict_9_4 = _T_15137 & _T_15138; // @[LoadQueue.scala 152:68:@15676.4]
  assign _T_15140 = entriesToCheck_9_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15678.4]
  assign _T_15141 = _T_15140 & addrKnown_9; // @[LoadQueue.scala 152:41:@15679.4]
  assign _T_15142 = addrQ_9 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15680.4]
  assign conflict_9_5 = _T_15141 & _T_15142; // @[LoadQueue.scala 152:68:@15681.4]
  assign _T_15144 = entriesToCheck_9_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15683.4]
  assign _T_15145 = _T_15144 & addrKnown_9; // @[LoadQueue.scala 152:41:@15684.4]
  assign _T_15146 = addrQ_9 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15685.4]
  assign conflict_9_6 = _T_15145 & _T_15146; // @[LoadQueue.scala 152:68:@15686.4]
  assign _T_15148 = entriesToCheck_9_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15688.4]
  assign _T_15149 = _T_15148 & addrKnown_9; // @[LoadQueue.scala 152:41:@15689.4]
  assign _T_15150 = addrQ_9 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15690.4]
  assign conflict_9_7 = _T_15149 & _T_15150; // @[LoadQueue.scala 152:68:@15691.4]
  assign _T_15152 = entriesToCheck_9_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15693.4]
  assign _T_15153 = _T_15152 & addrKnown_9; // @[LoadQueue.scala 152:41:@15694.4]
  assign _T_15154 = addrQ_9 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15695.4]
  assign conflict_9_8 = _T_15153 & _T_15154; // @[LoadQueue.scala 152:68:@15696.4]
  assign _T_15156 = entriesToCheck_9_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15698.4]
  assign _T_15157 = _T_15156 & addrKnown_9; // @[LoadQueue.scala 152:41:@15699.4]
  assign _T_15158 = addrQ_9 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15700.4]
  assign conflict_9_9 = _T_15157 & _T_15158; // @[LoadQueue.scala 152:68:@15701.4]
  assign _T_15160 = entriesToCheck_9_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15703.4]
  assign _T_15161 = _T_15160 & addrKnown_9; // @[LoadQueue.scala 152:41:@15704.4]
  assign _T_15162 = addrQ_9 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15705.4]
  assign conflict_9_10 = _T_15161 & _T_15162; // @[LoadQueue.scala 152:68:@15706.4]
  assign _T_15164 = entriesToCheck_9_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15708.4]
  assign _T_15165 = _T_15164 & addrKnown_9; // @[LoadQueue.scala 152:41:@15709.4]
  assign _T_15166 = addrQ_9 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15710.4]
  assign conflict_9_11 = _T_15165 & _T_15166; // @[LoadQueue.scala 152:68:@15711.4]
  assign _T_15168 = entriesToCheck_9_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15713.4]
  assign _T_15169 = _T_15168 & addrKnown_9; // @[LoadQueue.scala 152:41:@15714.4]
  assign _T_15170 = addrQ_9 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15715.4]
  assign conflict_9_12 = _T_15169 & _T_15170; // @[LoadQueue.scala 152:68:@15716.4]
  assign _T_15172 = entriesToCheck_9_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15718.4]
  assign _T_15173 = _T_15172 & addrKnown_9; // @[LoadQueue.scala 152:41:@15719.4]
  assign _T_15174 = addrQ_9 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15720.4]
  assign conflict_9_13 = _T_15173 & _T_15174; // @[LoadQueue.scala 152:68:@15721.4]
  assign _T_15176 = entriesToCheck_9_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15723.4]
  assign _T_15177 = _T_15176 & addrKnown_9; // @[LoadQueue.scala 152:41:@15724.4]
  assign _T_15178 = addrQ_9 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15725.4]
  assign conflict_9_14 = _T_15177 & _T_15178; // @[LoadQueue.scala 152:68:@15726.4]
  assign _T_15180 = entriesToCheck_9_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15728.4]
  assign _T_15181 = _T_15180 & addrKnown_9; // @[LoadQueue.scala 152:41:@15729.4]
  assign _T_15182 = addrQ_9 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15730.4]
  assign conflict_9_15 = _T_15181 & _T_15182; // @[LoadQueue.scala 152:68:@15731.4]
  assign _T_15184 = entriesToCheck_10_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15733.4]
  assign _T_15185 = _T_15184 & addrKnown_10; // @[LoadQueue.scala 152:41:@15734.4]
  assign _T_15186 = addrQ_10 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15735.4]
  assign conflict_10_0 = _T_15185 & _T_15186; // @[LoadQueue.scala 152:68:@15736.4]
  assign _T_15188 = entriesToCheck_10_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15738.4]
  assign _T_15189 = _T_15188 & addrKnown_10; // @[LoadQueue.scala 152:41:@15739.4]
  assign _T_15190 = addrQ_10 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15740.4]
  assign conflict_10_1 = _T_15189 & _T_15190; // @[LoadQueue.scala 152:68:@15741.4]
  assign _T_15192 = entriesToCheck_10_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15743.4]
  assign _T_15193 = _T_15192 & addrKnown_10; // @[LoadQueue.scala 152:41:@15744.4]
  assign _T_15194 = addrQ_10 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15745.4]
  assign conflict_10_2 = _T_15193 & _T_15194; // @[LoadQueue.scala 152:68:@15746.4]
  assign _T_15196 = entriesToCheck_10_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15748.4]
  assign _T_15197 = _T_15196 & addrKnown_10; // @[LoadQueue.scala 152:41:@15749.4]
  assign _T_15198 = addrQ_10 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15750.4]
  assign conflict_10_3 = _T_15197 & _T_15198; // @[LoadQueue.scala 152:68:@15751.4]
  assign _T_15200 = entriesToCheck_10_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15753.4]
  assign _T_15201 = _T_15200 & addrKnown_10; // @[LoadQueue.scala 152:41:@15754.4]
  assign _T_15202 = addrQ_10 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15755.4]
  assign conflict_10_4 = _T_15201 & _T_15202; // @[LoadQueue.scala 152:68:@15756.4]
  assign _T_15204 = entriesToCheck_10_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15758.4]
  assign _T_15205 = _T_15204 & addrKnown_10; // @[LoadQueue.scala 152:41:@15759.4]
  assign _T_15206 = addrQ_10 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15760.4]
  assign conflict_10_5 = _T_15205 & _T_15206; // @[LoadQueue.scala 152:68:@15761.4]
  assign _T_15208 = entriesToCheck_10_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15763.4]
  assign _T_15209 = _T_15208 & addrKnown_10; // @[LoadQueue.scala 152:41:@15764.4]
  assign _T_15210 = addrQ_10 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15765.4]
  assign conflict_10_6 = _T_15209 & _T_15210; // @[LoadQueue.scala 152:68:@15766.4]
  assign _T_15212 = entriesToCheck_10_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15768.4]
  assign _T_15213 = _T_15212 & addrKnown_10; // @[LoadQueue.scala 152:41:@15769.4]
  assign _T_15214 = addrQ_10 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15770.4]
  assign conflict_10_7 = _T_15213 & _T_15214; // @[LoadQueue.scala 152:68:@15771.4]
  assign _T_15216 = entriesToCheck_10_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15773.4]
  assign _T_15217 = _T_15216 & addrKnown_10; // @[LoadQueue.scala 152:41:@15774.4]
  assign _T_15218 = addrQ_10 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15775.4]
  assign conflict_10_8 = _T_15217 & _T_15218; // @[LoadQueue.scala 152:68:@15776.4]
  assign _T_15220 = entriesToCheck_10_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15778.4]
  assign _T_15221 = _T_15220 & addrKnown_10; // @[LoadQueue.scala 152:41:@15779.4]
  assign _T_15222 = addrQ_10 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15780.4]
  assign conflict_10_9 = _T_15221 & _T_15222; // @[LoadQueue.scala 152:68:@15781.4]
  assign _T_15224 = entriesToCheck_10_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15783.4]
  assign _T_15225 = _T_15224 & addrKnown_10; // @[LoadQueue.scala 152:41:@15784.4]
  assign _T_15226 = addrQ_10 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15785.4]
  assign conflict_10_10 = _T_15225 & _T_15226; // @[LoadQueue.scala 152:68:@15786.4]
  assign _T_15228 = entriesToCheck_10_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15788.4]
  assign _T_15229 = _T_15228 & addrKnown_10; // @[LoadQueue.scala 152:41:@15789.4]
  assign _T_15230 = addrQ_10 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15790.4]
  assign conflict_10_11 = _T_15229 & _T_15230; // @[LoadQueue.scala 152:68:@15791.4]
  assign _T_15232 = entriesToCheck_10_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15793.4]
  assign _T_15233 = _T_15232 & addrKnown_10; // @[LoadQueue.scala 152:41:@15794.4]
  assign _T_15234 = addrQ_10 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15795.4]
  assign conflict_10_12 = _T_15233 & _T_15234; // @[LoadQueue.scala 152:68:@15796.4]
  assign _T_15236 = entriesToCheck_10_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15798.4]
  assign _T_15237 = _T_15236 & addrKnown_10; // @[LoadQueue.scala 152:41:@15799.4]
  assign _T_15238 = addrQ_10 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15800.4]
  assign conflict_10_13 = _T_15237 & _T_15238; // @[LoadQueue.scala 152:68:@15801.4]
  assign _T_15240 = entriesToCheck_10_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15803.4]
  assign _T_15241 = _T_15240 & addrKnown_10; // @[LoadQueue.scala 152:41:@15804.4]
  assign _T_15242 = addrQ_10 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15805.4]
  assign conflict_10_14 = _T_15241 & _T_15242; // @[LoadQueue.scala 152:68:@15806.4]
  assign _T_15244 = entriesToCheck_10_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15808.4]
  assign _T_15245 = _T_15244 & addrKnown_10; // @[LoadQueue.scala 152:41:@15809.4]
  assign _T_15246 = addrQ_10 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15810.4]
  assign conflict_10_15 = _T_15245 & _T_15246; // @[LoadQueue.scala 152:68:@15811.4]
  assign _T_15248 = entriesToCheck_11_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15813.4]
  assign _T_15249 = _T_15248 & addrKnown_11; // @[LoadQueue.scala 152:41:@15814.4]
  assign _T_15250 = addrQ_11 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15815.4]
  assign conflict_11_0 = _T_15249 & _T_15250; // @[LoadQueue.scala 152:68:@15816.4]
  assign _T_15252 = entriesToCheck_11_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15818.4]
  assign _T_15253 = _T_15252 & addrKnown_11; // @[LoadQueue.scala 152:41:@15819.4]
  assign _T_15254 = addrQ_11 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15820.4]
  assign conflict_11_1 = _T_15253 & _T_15254; // @[LoadQueue.scala 152:68:@15821.4]
  assign _T_15256 = entriesToCheck_11_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15823.4]
  assign _T_15257 = _T_15256 & addrKnown_11; // @[LoadQueue.scala 152:41:@15824.4]
  assign _T_15258 = addrQ_11 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15825.4]
  assign conflict_11_2 = _T_15257 & _T_15258; // @[LoadQueue.scala 152:68:@15826.4]
  assign _T_15260 = entriesToCheck_11_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15828.4]
  assign _T_15261 = _T_15260 & addrKnown_11; // @[LoadQueue.scala 152:41:@15829.4]
  assign _T_15262 = addrQ_11 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15830.4]
  assign conflict_11_3 = _T_15261 & _T_15262; // @[LoadQueue.scala 152:68:@15831.4]
  assign _T_15264 = entriesToCheck_11_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15833.4]
  assign _T_15265 = _T_15264 & addrKnown_11; // @[LoadQueue.scala 152:41:@15834.4]
  assign _T_15266 = addrQ_11 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15835.4]
  assign conflict_11_4 = _T_15265 & _T_15266; // @[LoadQueue.scala 152:68:@15836.4]
  assign _T_15268 = entriesToCheck_11_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15838.4]
  assign _T_15269 = _T_15268 & addrKnown_11; // @[LoadQueue.scala 152:41:@15839.4]
  assign _T_15270 = addrQ_11 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15840.4]
  assign conflict_11_5 = _T_15269 & _T_15270; // @[LoadQueue.scala 152:68:@15841.4]
  assign _T_15272 = entriesToCheck_11_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15843.4]
  assign _T_15273 = _T_15272 & addrKnown_11; // @[LoadQueue.scala 152:41:@15844.4]
  assign _T_15274 = addrQ_11 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15845.4]
  assign conflict_11_6 = _T_15273 & _T_15274; // @[LoadQueue.scala 152:68:@15846.4]
  assign _T_15276 = entriesToCheck_11_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15848.4]
  assign _T_15277 = _T_15276 & addrKnown_11; // @[LoadQueue.scala 152:41:@15849.4]
  assign _T_15278 = addrQ_11 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15850.4]
  assign conflict_11_7 = _T_15277 & _T_15278; // @[LoadQueue.scala 152:68:@15851.4]
  assign _T_15280 = entriesToCheck_11_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15853.4]
  assign _T_15281 = _T_15280 & addrKnown_11; // @[LoadQueue.scala 152:41:@15854.4]
  assign _T_15282 = addrQ_11 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15855.4]
  assign conflict_11_8 = _T_15281 & _T_15282; // @[LoadQueue.scala 152:68:@15856.4]
  assign _T_15284 = entriesToCheck_11_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15858.4]
  assign _T_15285 = _T_15284 & addrKnown_11; // @[LoadQueue.scala 152:41:@15859.4]
  assign _T_15286 = addrQ_11 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15860.4]
  assign conflict_11_9 = _T_15285 & _T_15286; // @[LoadQueue.scala 152:68:@15861.4]
  assign _T_15288 = entriesToCheck_11_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15863.4]
  assign _T_15289 = _T_15288 & addrKnown_11; // @[LoadQueue.scala 152:41:@15864.4]
  assign _T_15290 = addrQ_11 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15865.4]
  assign conflict_11_10 = _T_15289 & _T_15290; // @[LoadQueue.scala 152:68:@15866.4]
  assign _T_15292 = entriesToCheck_11_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15868.4]
  assign _T_15293 = _T_15292 & addrKnown_11; // @[LoadQueue.scala 152:41:@15869.4]
  assign _T_15294 = addrQ_11 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15870.4]
  assign conflict_11_11 = _T_15293 & _T_15294; // @[LoadQueue.scala 152:68:@15871.4]
  assign _T_15296 = entriesToCheck_11_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15873.4]
  assign _T_15297 = _T_15296 & addrKnown_11; // @[LoadQueue.scala 152:41:@15874.4]
  assign _T_15298 = addrQ_11 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15875.4]
  assign conflict_11_12 = _T_15297 & _T_15298; // @[LoadQueue.scala 152:68:@15876.4]
  assign _T_15300 = entriesToCheck_11_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15878.4]
  assign _T_15301 = _T_15300 & addrKnown_11; // @[LoadQueue.scala 152:41:@15879.4]
  assign _T_15302 = addrQ_11 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15880.4]
  assign conflict_11_13 = _T_15301 & _T_15302; // @[LoadQueue.scala 152:68:@15881.4]
  assign _T_15304 = entriesToCheck_11_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15883.4]
  assign _T_15305 = _T_15304 & addrKnown_11; // @[LoadQueue.scala 152:41:@15884.4]
  assign _T_15306 = addrQ_11 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15885.4]
  assign conflict_11_14 = _T_15305 & _T_15306; // @[LoadQueue.scala 152:68:@15886.4]
  assign _T_15308 = entriesToCheck_11_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15888.4]
  assign _T_15309 = _T_15308 & addrKnown_11; // @[LoadQueue.scala 152:41:@15889.4]
  assign _T_15310 = addrQ_11 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15890.4]
  assign conflict_11_15 = _T_15309 & _T_15310; // @[LoadQueue.scala 152:68:@15891.4]
  assign _T_15312 = entriesToCheck_12_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15893.4]
  assign _T_15313 = _T_15312 & addrKnown_12; // @[LoadQueue.scala 152:41:@15894.4]
  assign _T_15314 = addrQ_12 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15895.4]
  assign conflict_12_0 = _T_15313 & _T_15314; // @[LoadQueue.scala 152:68:@15896.4]
  assign _T_15316 = entriesToCheck_12_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15898.4]
  assign _T_15317 = _T_15316 & addrKnown_12; // @[LoadQueue.scala 152:41:@15899.4]
  assign _T_15318 = addrQ_12 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15900.4]
  assign conflict_12_1 = _T_15317 & _T_15318; // @[LoadQueue.scala 152:68:@15901.4]
  assign _T_15320 = entriesToCheck_12_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15903.4]
  assign _T_15321 = _T_15320 & addrKnown_12; // @[LoadQueue.scala 152:41:@15904.4]
  assign _T_15322 = addrQ_12 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15905.4]
  assign conflict_12_2 = _T_15321 & _T_15322; // @[LoadQueue.scala 152:68:@15906.4]
  assign _T_15324 = entriesToCheck_12_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15908.4]
  assign _T_15325 = _T_15324 & addrKnown_12; // @[LoadQueue.scala 152:41:@15909.4]
  assign _T_15326 = addrQ_12 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15910.4]
  assign conflict_12_3 = _T_15325 & _T_15326; // @[LoadQueue.scala 152:68:@15911.4]
  assign _T_15328 = entriesToCheck_12_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15913.4]
  assign _T_15329 = _T_15328 & addrKnown_12; // @[LoadQueue.scala 152:41:@15914.4]
  assign _T_15330 = addrQ_12 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15915.4]
  assign conflict_12_4 = _T_15329 & _T_15330; // @[LoadQueue.scala 152:68:@15916.4]
  assign _T_15332 = entriesToCheck_12_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15918.4]
  assign _T_15333 = _T_15332 & addrKnown_12; // @[LoadQueue.scala 152:41:@15919.4]
  assign _T_15334 = addrQ_12 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@15920.4]
  assign conflict_12_5 = _T_15333 & _T_15334; // @[LoadQueue.scala 152:68:@15921.4]
  assign _T_15336 = entriesToCheck_12_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@15923.4]
  assign _T_15337 = _T_15336 & addrKnown_12; // @[LoadQueue.scala 152:41:@15924.4]
  assign _T_15338 = addrQ_12 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@15925.4]
  assign conflict_12_6 = _T_15337 & _T_15338; // @[LoadQueue.scala 152:68:@15926.4]
  assign _T_15340 = entriesToCheck_12_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@15928.4]
  assign _T_15341 = _T_15340 & addrKnown_12; // @[LoadQueue.scala 152:41:@15929.4]
  assign _T_15342 = addrQ_12 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@15930.4]
  assign conflict_12_7 = _T_15341 & _T_15342; // @[LoadQueue.scala 152:68:@15931.4]
  assign _T_15344 = entriesToCheck_12_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@15933.4]
  assign _T_15345 = _T_15344 & addrKnown_12; // @[LoadQueue.scala 152:41:@15934.4]
  assign _T_15346 = addrQ_12 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@15935.4]
  assign conflict_12_8 = _T_15345 & _T_15346; // @[LoadQueue.scala 152:68:@15936.4]
  assign _T_15348 = entriesToCheck_12_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@15938.4]
  assign _T_15349 = _T_15348 & addrKnown_12; // @[LoadQueue.scala 152:41:@15939.4]
  assign _T_15350 = addrQ_12 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@15940.4]
  assign conflict_12_9 = _T_15349 & _T_15350; // @[LoadQueue.scala 152:68:@15941.4]
  assign _T_15352 = entriesToCheck_12_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@15943.4]
  assign _T_15353 = _T_15352 & addrKnown_12; // @[LoadQueue.scala 152:41:@15944.4]
  assign _T_15354 = addrQ_12 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@15945.4]
  assign conflict_12_10 = _T_15353 & _T_15354; // @[LoadQueue.scala 152:68:@15946.4]
  assign _T_15356 = entriesToCheck_12_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@15948.4]
  assign _T_15357 = _T_15356 & addrKnown_12; // @[LoadQueue.scala 152:41:@15949.4]
  assign _T_15358 = addrQ_12 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@15950.4]
  assign conflict_12_11 = _T_15357 & _T_15358; // @[LoadQueue.scala 152:68:@15951.4]
  assign _T_15360 = entriesToCheck_12_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@15953.4]
  assign _T_15361 = _T_15360 & addrKnown_12; // @[LoadQueue.scala 152:41:@15954.4]
  assign _T_15362 = addrQ_12 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@15955.4]
  assign conflict_12_12 = _T_15361 & _T_15362; // @[LoadQueue.scala 152:68:@15956.4]
  assign _T_15364 = entriesToCheck_12_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@15958.4]
  assign _T_15365 = _T_15364 & addrKnown_12; // @[LoadQueue.scala 152:41:@15959.4]
  assign _T_15366 = addrQ_12 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@15960.4]
  assign conflict_12_13 = _T_15365 & _T_15366; // @[LoadQueue.scala 152:68:@15961.4]
  assign _T_15368 = entriesToCheck_12_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@15963.4]
  assign _T_15369 = _T_15368 & addrKnown_12; // @[LoadQueue.scala 152:41:@15964.4]
  assign _T_15370 = addrQ_12 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@15965.4]
  assign conflict_12_14 = _T_15369 & _T_15370; // @[LoadQueue.scala 152:68:@15966.4]
  assign _T_15372 = entriesToCheck_12_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@15968.4]
  assign _T_15373 = _T_15372 & addrKnown_12; // @[LoadQueue.scala 152:41:@15969.4]
  assign _T_15374 = addrQ_12 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@15970.4]
  assign conflict_12_15 = _T_15373 & _T_15374; // @[LoadQueue.scala 152:68:@15971.4]
  assign _T_15376 = entriesToCheck_13_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@15973.4]
  assign _T_15377 = _T_15376 & addrKnown_13; // @[LoadQueue.scala 152:41:@15974.4]
  assign _T_15378 = addrQ_13 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@15975.4]
  assign conflict_13_0 = _T_15377 & _T_15378; // @[LoadQueue.scala 152:68:@15976.4]
  assign _T_15380 = entriesToCheck_13_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@15978.4]
  assign _T_15381 = _T_15380 & addrKnown_13; // @[LoadQueue.scala 152:41:@15979.4]
  assign _T_15382 = addrQ_13 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@15980.4]
  assign conflict_13_1 = _T_15381 & _T_15382; // @[LoadQueue.scala 152:68:@15981.4]
  assign _T_15384 = entriesToCheck_13_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@15983.4]
  assign _T_15385 = _T_15384 & addrKnown_13; // @[LoadQueue.scala 152:41:@15984.4]
  assign _T_15386 = addrQ_13 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@15985.4]
  assign conflict_13_2 = _T_15385 & _T_15386; // @[LoadQueue.scala 152:68:@15986.4]
  assign _T_15388 = entriesToCheck_13_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@15988.4]
  assign _T_15389 = _T_15388 & addrKnown_13; // @[LoadQueue.scala 152:41:@15989.4]
  assign _T_15390 = addrQ_13 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@15990.4]
  assign conflict_13_3 = _T_15389 & _T_15390; // @[LoadQueue.scala 152:68:@15991.4]
  assign _T_15392 = entriesToCheck_13_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@15993.4]
  assign _T_15393 = _T_15392 & addrKnown_13; // @[LoadQueue.scala 152:41:@15994.4]
  assign _T_15394 = addrQ_13 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@15995.4]
  assign conflict_13_4 = _T_15393 & _T_15394; // @[LoadQueue.scala 152:68:@15996.4]
  assign _T_15396 = entriesToCheck_13_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@15998.4]
  assign _T_15397 = _T_15396 & addrKnown_13; // @[LoadQueue.scala 152:41:@15999.4]
  assign _T_15398 = addrQ_13 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@16000.4]
  assign conflict_13_5 = _T_15397 & _T_15398; // @[LoadQueue.scala 152:68:@16001.4]
  assign _T_15400 = entriesToCheck_13_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@16003.4]
  assign _T_15401 = _T_15400 & addrKnown_13; // @[LoadQueue.scala 152:41:@16004.4]
  assign _T_15402 = addrQ_13 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@16005.4]
  assign conflict_13_6 = _T_15401 & _T_15402; // @[LoadQueue.scala 152:68:@16006.4]
  assign _T_15404 = entriesToCheck_13_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@16008.4]
  assign _T_15405 = _T_15404 & addrKnown_13; // @[LoadQueue.scala 152:41:@16009.4]
  assign _T_15406 = addrQ_13 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@16010.4]
  assign conflict_13_7 = _T_15405 & _T_15406; // @[LoadQueue.scala 152:68:@16011.4]
  assign _T_15408 = entriesToCheck_13_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@16013.4]
  assign _T_15409 = _T_15408 & addrKnown_13; // @[LoadQueue.scala 152:41:@16014.4]
  assign _T_15410 = addrQ_13 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@16015.4]
  assign conflict_13_8 = _T_15409 & _T_15410; // @[LoadQueue.scala 152:68:@16016.4]
  assign _T_15412 = entriesToCheck_13_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@16018.4]
  assign _T_15413 = _T_15412 & addrKnown_13; // @[LoadQueue.scala 152:41:@16019.4]
  assign _T_15414 = addrQ_13 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@16020.4]
  assign conflict_13_9 = _T_15413 & _T_15414; // @[LoadQueue.scala 152:68:@16021.4]
  assign _T_15416 = entriesToCheck_13_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@16023.4]
  assign _T_15417 = _T_15416 & addrKnown_13; // @[LoadQueue.scala 152:41:@16024.4]
  assign _T_15418 = addrQ_13 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@16025.4]
  assign conflict_13_10 = _T_15417 & _T_15418; // @[LoadQueue.scala 152:68:@16026.4]
  assign _T_15420 = entriesToCheck_13_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@16028.4]
  assign _T_15421 = _T_15420 & addrKnown_13; // @[LoadQueue.scala 152:41:@16029.4]
  assign _T_15422 = addrQ_13 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@16030.4]
  assign conflict_13_11 = _T_15421 & _T_15422; // @[LoadQueue.scala 152:68:@16031.4]
  assign _T_15424 = entriesToCheck_13_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@16033.4]
  assign _T_15425 = _T_15424 & addrKnown_13; // @[LoadQueue.scala 152:41:@16034.4]
  assign _T_15426 = addrQ_13 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@16035.4]
  assign conflict_13_12 = _T_15425 & _T_15426; // @[LoadQueue.scala 152:68:@16036.4]
  assign _T_15428 = entriesToCheck_13_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@16038.4]
  assign _T_15429 = _T_15428 & addrKnown_13; // @[LoadQueue.scala 152:41:@16039.4]
  assign _T_15430 = addrQ_13 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@16040.4]
  assign conflict_13_13 = _T_15429 & _T_15430; // @[LoadQueue.scala 152:68:@16041.4]
  assign _T_15432 = entriesToCheck_13_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@16043.4]
  assign _T_15433 = _T_15432 & addrKnown_13; // @[LoadQueue.scala 152:41:@16044.4]
  assign _T_15434 = addrQ_13 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@16045.4]
  assign conflict_13_14 = _T_15433 & _T_15434; // @[LoadQueue.scala 152:68:@16046.4]
  assign _T_15436 = entriesToCheck_13_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@16048.4]
  assign _T_15437 = _T_15436 & addrKnown_13; // @[LoadQueue.scala 152:41:@16049.4]
  assign _T_15438 = addrQ_13 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@16050.4]
  assign conflict_13_15 = _T_15437 & _T_15438; // @[LoadQueue.scala 152:68:@16051.4]
  assign _T_15440 = entriesToCheck_14_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@16053.4]
  assign _T_15441 = _T_15440 & addrKnown_14; // @[LoadQueue.scala 152:41:@16054.4]
  assign _T_15442 = addrQ_14 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@16055.4]
  assign conflict_14_0 = _T_15441 & _T_15442; // @[LoadQueue.scala 152:68:@16056.4]
  assign _T_15444 = entriesToCheck_14_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@16058.4]
  assign _T_15445 = _T_15444 & addrKnown_14; // @[LoadQueue.scala 152:41:@16059.4]
  assign _T_15446 = addrQ_14 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@16060.4]
  assign conflict_14_1 = _T_15445 & _T_15446; // @[LoadQueue.scala 152:68:@16061.4]
  assign _T_15448 = entriesToCheck_14_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@16063.4]
  assign _T_15449 = _T_15448 & addrKnown_14; // @[LoadQueue.scala 152:41:@16064.4]
  assign _T_15450 = addrQ_14 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@16065.4]
  assign conflict_14_2 = _T_15449 & _T_15450; // @[LoadQueue.scala 152:68:@16066.4]
  assign _T_15452 = entriesToCheck_14_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@16068.4]
  assign _T_15453 = _T_15452 & addrKnown_14; // @[LoadQueue.scala 152:41:@16069.4]
  assign _T_15454 = addrQ_14 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@16070.4]
  assign conflict_14_3 = _T_15453 & _T_15454; // @[LoadQueue.scala 152:68:@16071.4]
  assign _T_15456 = entriesToCheck_14_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@16073.4]
  assign _T_15457 = _T_15456 & addrKnown_14; // @[LoadQueue.scala 152:41:@16074.4]
  assign _T_15458 = addrQ_14 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@16075.4]
  assign conflict_14_4 = _T_15457 & _T_15458; // @[LoadQueue.scala 152:68:@16076.4]
  assign _T_15460 = entriesToCheck_14_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@16078.4]
  assign _T_15461 = _T_15460 & addrKnown_14; // @[LoadQueue.scala 152:41:@16079.4]
  assign _T_15462 = addrQ_14 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@16080.4]
  assign conflict_14_5 = _T_15461 & _T_15462; // @[LoadQueue.scala 152:68:@16081.4]
  assign _T_15464 = entriesToCheck_14_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@16083.4]
  assign _T_15465 = _T_15464 & addrKnown_14; // @[LoadQueue.scala 152:41:@16084.4]
  assign _T_15466 = addrQ_14 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@16085.4]
  assign conflict_14_6 = _T_15465 & _T_15466; // @[LoadQueue.scala 152:68:@16086.4]
  assign _T_15468 = entriesToCheck_14_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@16088.4]
  assign _T_15469 = _T_15468 & addrKnown_14; // @[LoadQueue.scala 152:41:@16089.4]
  assign _T_15470 = addrQ_14 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@16090.4]
  assign conflict_14_7 = _T_15469 & _T_15470; // @[LoadQueue.scala 152:68:@16091.4]
  assign _T_15472 = entriesToCheck_14_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@16093.4]
  assign _T_15473 = _T_15472 & addrKnown_14; // @[LoadQueue.scala 152:41:@16094.4]
  assign _T_15474 = addrQ_14 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@16095.4]
  assign conflict_14_8 = _T_15473 & _T_15474; // @[LoadQueue.scala 152:68:@16096.4]
  assign _T_15476 = entriesToCheck_14_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@16098.4]
  assign _T_15477 = _T_15476 & addrKnown_14; // @[LoadQueue.scala 152:41:@16099.4]
  assign _T_15478 = addrQ_14 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@16100.4]
  assign conflict_14_9 = _T_15477 & _T_15478; // @[LoadQueue.scala 152:68:@16101.4]
  assign _T_15480 = entriesToCheck_14_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@16103.4]
  assign _T_15481 = _T_15480 & addrKnown_14; // @[LoadQueue.scala 152:41:@16104.4]
  assign _T_15482 = addrQ_14 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@16105.4]
  assign conflict_14_10 = _T_15481 & _T_15482; // @[LoadQueue.scala 152:68:@16106.4]
  assign _T_15484 = entriesToCheck_14_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@16108.4]
  assign _T_15485 = _T_15484 & addrKnown_14; // @[LoadQueue.scala 152:41:@16109.4]
  assign _T_15486 = addrQ_14 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@16110.4]
  assign conflict_14_11 = _T_15485 & _T_15486; // @[LoadQueue.scala 152:68:@16111.4]
  assign _T_15488 = entriesToCheck_14_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@16113.4]
  assign _T_15489 = _T_15488 & addrKnown_14; // @[LoadQueue.scala 152:41:@16114.4]
  assign _T_15490 = addrQ_14 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@16115.4]
  assign conflict_14_12 = _T_15489 & _T_15490; // @[LoadQueue.scala 152:68:@16116.4]
  assign _T_15492 = entriesToCheck_14_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@16118.4]
  assign _T_15493 = _T_15492 & addrKnown_14; // @[LoadQueue.scala 152:41:@16119.4]
  assign _T_15494 = addrQ_14 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@16120.4]
  assign conflict_14_13 = _T_15493 & _T_15494; // @[LoadQueue.scala 152:68:@16121.4]
  assign _T_15496 = entriesToCheck_14_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@16123.4]
  assign _T_15497 = _T_15496 & addrKnown_14; // @[LoadQueue.scala 152:41:@16124.4]
  assign _T_15498 = addrQ_14 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@16125.4]
  assign conflict_14_14 = _T_15497 & _T_15498; // @[LoadQueue.scala 152:68:@16126.4]
  assign _T_15500 = entriesToCheck_14_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@16128.4]
  assign _T_15501 = _T_15500 & addrKnown_14; // @[LoadQueue.scala 152:41:@16129.4]
  assign _T_15502 = addrQ_14 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@16130.4]
  assign conflict_14_15 = _T_15501 & _T_15502; // @[LoadQueue.scala 152:68:@16131.4]
  assign _T_15504 = entriesToCheck_15_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@16133.4]
  assign _T_15505 = _T_15504 & addrKnown_15; // @[LoadQueue.scala 152:41:@16134.4]
  assign _T_15506 = addrQ_15 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@16135.4]
  assign conflict_15_0 = _T_15505 & _T_15506; // @[LoadQueue.scala 152:68:@16136.4]
  assign _T_15508 = entriesToCheck_15_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@16138.4]
  assign _T_15509 = _T_15508 & addrKnown_15; // @[LoadQueue.scala 152:41:@16139.4]
  assign _T_15510 = addrQ_15 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@16140.4]
  assign conflict_15_1 = _T_15509 & _T_15510; // @[LoadQueue.scala 152:68:@16141.4]
  assign _T_15512 = entriesToCheck_15_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@16143.4]
  assign _T_15513 = _T_15512 & addrKnown_15; // @[LoadQueue.scala 152:41:@16144.4]
  assign _T_15514 = addrQ_15 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@16145.4]
  assign conflict_15_2 = _T_15513 & _T_15514; // @[LoadQueue.scala 152:68:@16146.4]
  assign _T_15516 = entriesToCheck_15_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@16148.4]
  assign _T_15517 = _T_15516 & addrKnown_15; // @[LoadQueue.scala 152:41:@16149.4]
  assign _T_15518 = addrQ_15 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@16150.4]
  assign conflict_15_3 = _T_15517 & _T_15518; // @[LoadQueue.scala 152:68:@16151.4]
  assign _T_15520 = entriesToCheck_15_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@16153.4]
  assign _T_15521 = _T_15520 & addrKnown_15; // @[LoadQueue.scala 152:41:@16154.4]
  assign _T_15522 = addrQ_15 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@16155.4]
  assign conflict_15_4 = _T_15521 & _T_15522; // @[LoadQueue.scala 152:68:@16156.4]
  assign _T_15524 = entriesToCheck_15_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@16158.4]
  assign _T_15525 = _T_15524 & addrKnown_15; // @[LoadQueue.scala 152:41:@16159.4]
  assign _T_15526 = addrQ_15 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@16160.4]
  assign conflict_15_5 = _T_15525 & _T_15526; // @[LoadQueue.scala 152:68:@16161.4]
  assign _T_15528 = entriesToCheck_15_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@16163.4]
  assign _T_15529 = _T_15528 & addrKnown_15; // @[LoadQueue.scala 152:41:@16164.4]
  assign _T_15530 = addrQ_15 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@16165.4]
  assign conflict_15_6 = _T_15529 & _T_15530; // @[LoadQueue.scala 152:68:@16166.4]
  assign _T_15532 = entriesToCheck_15_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@16168.4]
  assign _T_15533 = _T_15532 & addrKnown_15; // @[LoadQueue.scala 152:41:@16169.4]
  assign _T_15534 = addrQ_15 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@16170.4]
  assign conflict_15_7 = _T_15533 & _T_15534; // @[LoadQueue.scala 152:68:@16171.4]
  assign _T_15536 = entriesToCheck_15_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@16173.4]
  assign _T_15537 = _T_15536 & addrKnown_15; // @[LoadQueue.scala 152:41:@16174.4]
  assign _T_15538 = addrQ_15 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@16175.4]
  assign conflict_15_8 = _T_15537 & _T_15538; // @[LoadQueue.scala 152:68:@16176.4]
  assign _T_15540 = entriesToCheck_15_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@16178.4]
  assign _T_15541 = _T_15540 & addrKnown_15; // @[LoadQueue.scala 152:41:@16179.4]
  assign _T_15542 = addrQ_15 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@16180.4]
  assign conflict_15_9 = _T_15541 & _T_15542; // @[LoadQueue.scala 152:68:@16181.4]
  assign _T_15544 = entriesToCheck_15_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@16183.4]
  assign _T_15545 = _T_15544 & addrKnown_15; // @[LoadQueue.scala 152:41:@16184.4]
  assign _T_15546 = addrQ_15 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@16185.4]
  assign conflict_15_10 = _T_15545 & _T_15546; // @[LoadQueue.scala 152:68:@16186.4]
  assign _T_15548 = entriesToCheck_15_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@16188.4]
  assign _T_15549 = _T_15548 & addrKnown_15; // @[LoadQueue.scala 152:41:@16189.4]
  assign _T_15550 = addrQ_15 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@16190.4]
  assign conflict_15_11 = _T_15549 & _T_15550; // @[LoadQueue.scala 152:68:@16191.4]
  assign _T_15552 = entriesToCheck_15_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@16193.4]
  assign _T_15553 = _T_15552 & addrKnown_15; // @[LoadQueue.scala 152:41:@16194.4]
  assign _T_15554 = addrQ_15 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@16195.4]
  assign conflict_15_12 = _T_15553 & _T_15554; // @[LoadQueue.scala 152:68:@16196.4]
  assign _T_15556 = entriesToCheck_15_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@16198.4]
  assign _T_15557 = _T_15556 & addrKnown_15; // @[LoadQueue.scala 152:41:@16199.4]
  assign _T_15558 = addrQ_15 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@16200.4]
  assign conflict_15_13 = _T_15557 & _T_15558; // @[LoadQueue.scala 152:68:@16201.4]
  assign _T_15560 = entriesToCheck_15_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@16203.4]
  assign _T_15561 = _T_15560 & addrKnown_15; // @[LoadQueue.scala 152:41:@16204.4]
  assign _T_15562 = addrQ_15 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@16205.4]
  assign conflict_15_14 = _T_15561 & _T_15562; // @[LoadQueue.scala 152:68:@16206.4]
  assign _T_15564 = entriesToCheck_15_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@16208.4]
  assign _T_15565 = _T_15564 & addrKnown_15; // @[LoadQueue.scala 152:41:@16209.4]
  assign _T_15566 = addrQ_15 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@16210.4]
  assign conflict_15_15 = _T_15565 & _T_15566; // @[LoadQueue.scala 152:68:@16211.4]
  assign _T_16799 = io_storeAddrDone_0 == 1'h0; // @[LoadQueue.scala 163:13:@16214.4]
  assign storeAddrNotKnownFlags_0_0 = _T_16799 & entriesToCheck_0_0; // @[LoadQueue.scala 163:19:@16215.4]
  assign _T_16802 = io_storeAddrDone_1 == 1'h0; // @[LoadQueue.scala 163:13:@16216.4]
  assign storeAddrNotKnownFlags_0_1 = _T_16802 & entriesToCheck_0_1; // @[LoadQueue.scala 163:19:@16217.4]
  assign _T_16805 = io_storeAddrDone_2 == 1'h0; // @[LoadQueue.scala 163:13:@16218.4]
  assign storeAddrNotKnownFlags_0_2 = _T_16805 & entriesToCheck_0_2; // @[LoadQueue.scala 163:19:@16219.4]
  assign _T_16808 = io_storeAddrDone_3 == 1'h0; // @[LoadQueue.scala 163:13:@16220.4]
  assign storeAddrNotKnownFlags_0_3 = _T_16808 & entriesToCheck_0_3; // @[LoadQueue.scala 163:19:@16221.4]
  assign _T_16811 = io_storeAddrDone_4 == 1'h0; // @[LoadQueue.scala 163:13:@16222.4]
  assign storeAddrNotKnownFlags_0_4 = _T_16811 & entriesToCheck_0_4; // @[LoadQueue.scala 163:19:@16223.4]
  assign _T_16814 = io_storeAddrDone_5 == 1'h0; // @[LoadQueue.scala 163:13:@16224.4]
  assign storeAddrNotKnownFlags_0_5 = _T_16814 & entriesToCheck_0_5; // @[LoadQueue.scala 163:19:@16225.4]
  assign _T_16817 = io_storeAddrDone_6 == 1'h0; // @[LoadQueue.scala 163:13:@16226.4]
  assign storeAddrNotKnownFlags_0_6 = _T_16817 & entriesToCheck_0_6; // @[LoadQueue.scala 163:19:@16227.4]
  assign _T_16820 = io_storeAddrDone_7 == 1'h0; // @[LoadQueue.scala 163:13:@16228.4]
  assign storeAddrNotKnownFlags_0_7 = _T_16820 & entriesToCheck_0_7; // @[LoadQueue.scala 163:19:@16229.4]
  assign _T_16823 = io_storeAddrDone_8 == 1'h0; // @[LoadQueue.scala 163:13:@16230.4]
  assign storeAddrNotKnownFlags_0_8 = _T_16823 & entriesToCheck_0_8; // @[LoadQueue.scala 163:19:@16231.4]
  assign _T_16826 = io_storeAddrDone_9 == 1'h0; // @[LoadQueue.scala 163:13:@16232.4]
  assign storeAddrNotKnownFlags_0_9 = _T_16826 & entriesToCheck_0_9; // @[LoadQueue.scala 163:19:@16233.4]
  assign _T_16829 = io_storeAddrDone_10 == 1'h0; // @[LoadQueue.scala 163:13:@16234.4]
  assign storeAddrNotKnownFlags_0_10 = _T_16829 & entriesToCheck_0_10; // @[LoadQueue.scala 163:19:@16235.4]
  assign _T_16832 = io_storeAddrDone_11 == 1'h0; // @[LoadQueue.scala 163:13:@16236.4]
  assign storeAddrNotKnownFlags_0_11 = _T_16832 & entriesToCheck_0_11; // @[LoadQueue.scala 163:19:@16237.4]
  assign _T_16835 = io_storeAddrDone_12 == 1'h0; // @[LoadQueue.scala 163:13:@16238.4]
  assign storeAddrNotKnownFlags_0_12 = _T_16835 & entriesToCheck_0_12; // @[LoadQueue.scala 163:19:@16239.4]
  assign _T_16838 = io_storeAddrDone_13 == 1'h0; // @[LoadQueue.scala 163:13:@16240.4]
  assign storeAddrNotKnownFlags_0_13 = _T_16838 & entriesToCheck_0_13; // @[LoadQueue.scala 163:19:@16241.4]
  assign _T_16841 = io_storeAddrDone_14 == 1'h0; // @[LoadQueue.scala 163:13:@16242.4]
  assign storeAddrNotKnownFlags_0_14 = _T_16841 & entriesToCheck_0_14; // @[LoadQueue.scala 163:19:@16243.4]
  assign _T_16844 = io_storeAddrDone_15 == 1'h0; // @[LoadQueue.scala 163:13:@16244.4]
  assign storeAddrNotKnownFlags_0_15 = _T_16844 & entriesToCheck_0_15; // @[LoadQueue.scala 163:19:@16245.4]
  assign storeAddrNotKnownFlags_1_0 = _T_16799 & entriesToCheck_1_0; // @[LoadQueue.scala 163:19:@16263.4]
  assign storeAddrNotKnownFlags_1_1 = _T_16802 & entriesToCheck_1_1; // @[LoadQueue.scala 163:19:@16265.4]
  assign storeAddrNotKnownFlags_1_2 = _T_16805 & entriesToCheck_1_2; // @[LoadQueue.scala 163:19:@16267.4]
  assign storeAddrNotKnownFlags_1_3 = _T_16808 & entriesToCheck_1_3; // @[LoadQueue.scala 163:19:@16269.4]
  assign storeAddrNotKnownFlags_1_4 = _T_16811 & entriesToCheck_1_4; // @[LoadQueue.scala 163:19:@16271.4]
  assign storeAddrNotKnownFlags_1_5 = _T_16814 & entriesToCheck_1_5; // @[LoadQueue.scala 163:19:@16273.4]
  assign storeAddrNotKnownFlags_1_6 = _T_16817 & entriesToCheck_1_6; // @[LoadQueue.scala 163:19:@16275.4]
  assign storeAddrNotKnownFlags_1_7 = _T_16820 & entriesToCheck_1_7; // @[LoadQueue.scala 163:19:@16277.4]
  assign storeAddrNotKnownFlags_1_8 = _T_16823 & entriesToCheck_1_8; // @[LoadQueue.scala 163:19:@16279.4]
  assign storeAddrNotKnownFlags_1_9 = _T_16826 & entriesToCheck_1_9; // @[LoadQueue.scala 163:19:@16281.4]
  assign storeAddrNotKnownFlags_1_10 = _T_16829 & entriesToCheck_1_10; // @[LoadQueue.scala 163:19:@16283.4]
  assign storeAddrNotKnownFlags_1_11 = _T_16832 & entriesToCheck_1_11; // @[LoadQueue.scala 163:19:@16285.4]
  assign storeAddrNotKnownFlags_1_12 = _T_16835 & entriesToCheck_1_12; // @[LoadQueue.scala 163:19:@16287.4]
  assign storeAddrNotKnownFlags_1_13 = _T_16838 & entriesToCheck_1_13; // @[LoadQueue.scala 163:19:@16289.4]
  assign storeAddrNotKnownFlags_1_14 = _T_16841 & entriesToCheck_1_14; // @[LoadQueue.scala 163:19:@16291.4]
  assign storeAddrNotKnownFlags_1_15 = _T_16844 & entriesToCheck_1_15; // @[LoadQueue.scala 163:19:@16293.4]
  assign storeAddrNotKnownFlags_2_0 = _T_16799 & entriesToCheck_2_0; // @[LoadQueue.scala 163:19:@16311.4]
  assign storeAddrNotKnownFlags_2_1 = _T_16802 & entriesToCheck_2_1; // @[LoadQueue.scala 163:19:@16313.4]
  assign storeAddrNotKnownFlags_2_2 = _T_16805 & entriesToCheck_2_2; // @[LoadQueue.scala 163:19:@16315.4]
  assign storeAddrNotKnownFlags_2_3 = _T_16808 & entriesToCheck_2_3; // @[LoadQueue.scala 163:19:@16317.4]
  assign storeAddrNotKnownFlags_2_4 = _T_16811 & entriesToCheck_2_4; // @[LoadQueue.scala 163:19:@16319.4]
  assign storeAddrNotKnownFlags_2_5 = _T_16814 & entriesToCheck_2_5; // @[LoadQueue.scala 163:19:@16321.4]
  assign storeAddrNotKnownFlags_2_6 = _T_16817 & entriesToCheck_2_6; // @[LoadQueue.scala 163:19:@16323.4]
  assign storeAddrNotKnownFlags_2_7 = _T_16820 & entriesToCheck_2_7; // @[LoadQueue.scala 163:19:@16325.4]
  assign storeAddrNotKnownFlags_2_8 = _T_16823 & entriesToCheck_2_8; // @[LoadQueue.scala 163:19:@16327.4]
  assign storeAddrNotKnownFlags_2_9 = _T_16826 & entriesToCheck_2_9; // @[LoadQueue.scala 163:19:@16329.4]
  assign storeAddrNotKnownFlags_2_10 = _T_16829 & entriesToCheck_2_10; // @[LoadQueue.scala 163:19:@16331.4]
  assign storeAddrNotKnownFlags_2_11 = _T_16832 & entriesToCheck_2_11; // @[LoadQueue.scala 163:19:@16333.4]
  assign storeAddrNotKnownFlags_2_12 = _T_16835 & entriesToCheck_2_12; // @[LoadQueue.scala 163:19:@16335.4]
  assign storeAddrNotKnownFlags_2_13 = _T_16838 & entriesToCheck_2_13; // @[LoadQueue.scala 163:19:@16337.4]
  assign storeAddrNotKnownFlags_2_14 = _T_16841 & entriesToCheck_2_14; // @[LoadQueue.scala 163:19:@16339.4]
  assign storeAddrNotKnownFlags_2_15 = _T_16844 & entriesToCheck_2_15; // @[LoadQueue.scala 163:19:@16341.4]
  assign storeAddrNotKnownFlags_3_0 = _T_16799 & entriesToCheck_3_0; // @[LoadQueue.scala 163:19:@16359.4]
  assign storeAddrNotKnownFlags_3_1 = _T_16802 & entriesToCheck_3_1; // @[LoadQueue.scala 163:19:@16361.4]
  assign storeAddrNotKnownFlags_3_2 = _T_16805 & entriesToCheck_3_2; // @[LoadQueue.scala 163:19:@16363.4]
  assign storeAddrNotKnownFlags_3_3 = _T_16808 & entriesToCheck_3_3; // @[LoadQueue.scala 163:19:@16365.4]
  assign storeAddrNotKnownFlags_3_4 = _T_16811 & entriesToCheck_3_4; // @[LoadQueue.scala 163:19:@16367.4]
  assign storeAddrNotKnownFlags_3_5 = _T_16814 & entriesToCheck_3_5; // @[LoadQueue.scala 163:19:@16369.4]
  assign storeAddrNotKnownFlags_3_6 = _T_16817 & entriesToCheck_3_6; // @[LoadQueue.scala 163:19:@16371.4]
  assign storeAddrNotKnownFlags_3_7 = _T_16820 & entriesToCheck_3_7; // @[LoadQueue.scala 163:19:@16373.4]
  assign storeAddrNotKnownFlags_3_8 = _T_16823 & entriesToCheck_3_8; // @[LoadQueue.scala 163:19:@16375.4]
  assign storeAddrNotKnownFlags_3_9 = _T_16826 & entriesToCheck_3_9; // @[LoadQueue.scala 163:19:@16377.4]
  assign storeAddrNotKnownFlags_3_10 = _T_16829 & entriesToCheck_3_10; // @[LoadQueue.scala 163:19:@16379.4]
  assign storeAddrNotKnownFlags_3_11 = _T_16832 & entriesToCheck_3_11; // @[LoadQueue.scala 163:19:@16381.4]
  assign storeAddrNotKnownFlags_3_12 = _T_16835 & entriesToCheck_3_12; // @[LoadQueue.scala 163:19:@16383.4]
  assign storeAddrNotKnownFlags_3_13 = _T_16838 & entriesToCheck_3_13; // @[LoadQueue.scala 163:19:@16385.4]
  assign storeAddrNotKnownFlags_3_14 = _T_16841 & entriesToCheck_3_14; // @[LoadQueue.scala 163:19:@16387.4]
  assign storeAddrNotKnownFlags_3_15 = _T_16844 & entriesToCheck_3_15; // @[LoadQueue.scala 163:19:@16389.4]
  assign storeAddrNotKnownFlags_4_0 = _T_16799 & entriesToCheck_4_0; // @[LoadQueue.scala 163:19:@16407.4]
  assign storeAddrNotKnownFlags_4_1 = _T_16802 & entriesToCheck_4_1; // @[LoadQueue.scala 163:19:@16409.4]
  assign storeAddrNotKnownFlags_4_2 = _T_16805 & entriesToCheck_4_2; // @[LoadQueue.scala 163:19:@16411.4]
  assign storeAddrNotKnownFlags_4_3 = _T_16808 & entriesToCheck_4_3; // @[LoadQueue.scala 163:19:@16413.4]
  assign storeAddrNotKnownFlags_4_4 = _T_16811 & entriesToCheck_4_4; // @[LoadQueue.scala 163:19:@16415.4]
  assign storeAddrNotKnownFlags_4_5 = _T_16814 & entriesToCheck_4_5; // @[LoadQueue.scala 163:19:@16417.4]
  assign storeAddrNotKnownFlags_4_6 = _T_16817 & entriesToCheck_4_6; // @[LoadQueue.scala 163:19:@16419.4]
  assign storeAddrNotKnownFlags_4_7 = _T_16820 & entriesToCheck_4_7; // @[LoadQueue.scala 163:19:@16421.4]
  assign storeAddrNotKnownFlags_4_8 = _T_16823 & entriesToCheck_4_8; // @[LoadQueue.scala 163:19:@16423.4]
  assign storeAddrNotKnownFlags_4_9 = _T_16826 & entriesToCheck_4_9; // @[LoadQueue.scala 163:19:@16425.4]
  assign storeAddrNotKnownFlags_4_10 = _T_16829 & entriesToCheck_4_10; // @[LoadQueue.scala 163:19:@16427.4]
  assign storeAddrNotKnownFlags_4_11 = _T_16832 & entriesToCheck_4_11; // @[LoadQueue.scala 163:19:@16429.4]
  assign storeAddrNotKnownFlags_4_12 = _T_16835 & entriesToCheck_4_12; // @[LoadQueue.scala 163:19:@16431.4]
  assign storeAddrNotKnownFlags_4_13 = _T_16838 & entriesToCheck_4_13; // @[LoadQueue.scala 163:19:@16433.4]
  assign storeAddrNotKnownFlags_4_14 = _T_16841 & entriesToCheck_4_14; // @[LoadQueue.scala 163:19:@16435.4]
  assign storeAddrNotKnownFlags_4_15 = _T_16844 & entriesToCheck_4_15; // @[LoadQueue.scala 163:19:@16437.4]
  assign storeAddrNotKnownFlags_5_0 = _T_16799 & entriesToCheck_5_0; // @[LoadQueue.scala 163:19:@16455.4]
  assign storeAddrNotKnownFlags_5_1 = _T_16802 & entriesToCheck_5_1; // @[LoadQueue.scala 163:19:@16457.4]
  assign storeAddrNotKnownFlags_5_2 = _T_16805 & entriesToCheck_5_2; // @[LoadQueue.scala 163:19:@16459.4]
  assign storeAddrNotKnownFlags_5_3 = _T_16808 & entriesToCheck_5_3; // @[LoadQueue.scala 163:19:@16461.4]
  assign storeAddrNotKnownFlags_5_4 = _T_16811 & entriesToCheck_5_4; // @[LoadQueue.scala 163:19:@16463.4]
  assign storeAddrNotKnownFlags_5_5 = _T_16814 & entriesToCheck_5_5; // @[LoadQueue.scala 163:19:@16465.4]
  assign storeAddrNotKnownFlags_5_6 = _T_16817 & entriesToCheck_5_6; // @[LoadQueue.scala 163:19:@16467.4]
  assign storeAddrNotKnownFlags_5_7 = _T_16820 & entriesToCheck_5_7; // @[LoadQueue.scala 163:19:@16469.4]
  assign storeAddrNotKnownFlags_5_8 = _T_16823 & entriesToCheck_5_8; // @[LoadQueue.scala 163:19:@16471.4]
  assign storeAddrNotKnownFlags_5_9 = _T_16826 & entriesToCheck_5_9; // @[LoadQueue.scala 163:19:@16473.4]
  assign storeAddrNotKnownFlags_5_10 = _T_16829 & entriesToCheck_5_10; // @[LoadQueue.scala 163:19:@16475.4]
  assign storeAddrNotKnownFlags_5_11 = _T_16832 & entriesToCheck_5_11; // @[LoadQueue.scala 163:19:@16477.4]
  assign storeAddrNotKnownFlags_5_12 = _T_16835 & entriesToCheck_5_12; // @[LoadQueue.scala 163:19:@16479.4]
  assign storeAddrNotKnownFlags_5_13 = _T_16838 & entriesToCheck_5_13; // @[LoadQueue.scala 163:19:@16481.4]
  assign storeAddrNotKnownFlags_5_14 = _T_16841 & entriesToCheck_5_14; // @[LoadQueue.scala 163:19:@16483.4]
  assign storeAddrNotKnownFlags_5_15 = _T_16844 & entriesToCheck_5_15; // @[LoadQueue.scala 163:19:@16485.4]
  assign storeAddrNotKnownFlags_6_0 = _T_16799 & entriesToCheck_6_0; // @[LoadQueue.scala 163:19:@16503.4]
  assign storeAddrNotKnownFlags_6_1 = _T_16802 & entriesToCheck_6_1; // @[LoadQueue.scala 163:19:@16505.4]
  assign storeAddrNotKnownFlags_6_2 = _T_16805 & entriesToCheck_6_2; // @[LoadQueue.scala 163:19:@16507.4]
  assign storeAddrNotKnownFlags_6_3 = _T_16808 & entriesToCheck_6_3; // @[LoadQueue.scala 163:19:@16509.4]
  assign storeAddrNotKnownFlags_6_4 = _T_16811 & entriesToCheck_6_4; // @[LoadQueue.scala 163:19:@16511.4]
  assign storeAddrNotKnownFlags_6_5 = _T_16814 & entriesToCheck_6_5; // @[LoadQueue.scala 163:19:@16513.4]
  assign storeAddrNotKnownFlags_6_6 = _T_16817 & entriesToCheck_6_6; // @[LoadQueue.scala 163:19:@16515.4]
  assign storeAddrNotKnownFlags_6_7 = _T_16820 & entriesToCheck_6_7; // @[LoadQueue.scala 163:19:@16517.4]
  assign storeAddrNotKnownFlags_6_8 = _T_16823 & entriesToCheck_6_8; // @[LoadQueue.scala 163:19:@16519.4]
  assign storeAddrNotKnownFlags_6_9 = _T_16826 & entriesToCheck_6_9; // @[LoadQueue.scala 163:19:@16521.4]
  assign storeAddrNotKnownFlags_6_10 = _T_16829 & entriesToCheck_6_10; // @[LoadQueue.scala 163:19:@16523.4]
  assign storeAddrNotKnownFlags_6_11 = _T_16832 & entriesToCheck_6_11; // @[LoadQueue.scala 163:19:@16525.4]
  assign storeAddrNotKnownFlags_6_12 = _T_16835 & entriesToCheck_6_12; // @[LoadQueue.scala 163:19:@16527.4]
  assign storeAddrNotKnownFlags_6_13 = _T_16838 & entriesToCheck_6_13; // @[LoadQueue.scala 163:19:@16529.4]
  assign storeAddrNotKnownFlags_6_14 = _T_16841 & entriesToCheck_6_14; // @[LoadQueue.scala 163:19:@16531.4]
  assign storeAddrNotKnownFlags_6_15 = _T_16844 & entriesToCheck_6_15; // @[LoadQueue.scala 163:19:@16533.4]
  assign storeAddrNotKnownFlags_7_0 = _T_16799 & entriesToCheck_7_0; // @[LoadQueue.scala 163:19:@16551.4]
  assign storeAddrNotKnownFlags_7_1 = _T_16802 & entriesToCheck_7_1; // @[LoadQueue.scala 163:19:@16553.4]
  assign storeAddrNotKnownFlags_7_2 = _T_16805 & entriesToCheck_7_2; // @[LoadQueue.scala 163:19:@16555.4]
  assign storeAddrNotKnownFlags_7_3 = _T_16808 & entriesToCheck_7_3; // @[LoadQueue.scala 163:19:@16557.4]
  assign storeAddrNotKnownFlags_7_4 = _T_16811 & entriesToCheck_7_4; // @[LoadQueue.scala 163:19:@16559.4]
  assign storeAddrNotKnownFlags_7_5 = _T_16814 & entriesToCheck_7_5; // @[LoadQueue.scala 163:19:@16561.4]
  assign storeAddrNotKnownFlags_7_6 = _T_16817 & entriesToCheck_7_6; // @[LoadQueue.scala 163:19:@16563.4]
  assign storeAddrNotKnownFlags_7_7 = _T_16820 & entriesToCheck_7_7; // @[LoadQueue.scala 163:19:@16565.4]
  assign storeAddrNotKnownFlags_7_8 = _T_16823 & entriesToCheck_7_8; // @[LoadQueue.scala 163:19:@16567.4]
  assign storeAddrNotKnownFlags_7_9 = _T_16826 & entriesToCheck_7_9; // @[LoadQueue.scala 163:19:@16569.4]
  assign storeAddrNotKnownFlags_7_10 = _T_16829 & entriesToCheck_7_10; // @[LoadQueue.scala 163:19:@16571.4]
  assign storeAddrNotKnownFlags_7_11 = _T_16832 & entriesToCheck_7_11; // @[LoadQueue.scala 163:19:@16573.4]
  assign storeAddrNotKnownFlags_7_12 = _T_16835 & entriesToCheck_7_12; // @[LoadQueue.scala 163:19:@16575.4]
  assign storeAddrNotKnownFlags_7_13 = _T_16838 & entriesToCheck_7_13; // @[LoadQueue.scala 163:19:@16577.4]
  assign storeAddrNotKnownFlags_7_14 = _T_16841 & entriesToCheck_7_14; // @[LoadQueue.scala 163:19:@16579.4]
  assign storeAddrNotKnownFlags_7_15 = _T_16844 & entriesToCheck_7_15; // @[LoadQueue.scala 163:19:@16581.4]
  assign storeAddrNotKnownFlags_8_0 = _T_16799 & entriesToCheck_8_0; // @[LoadQueue.scala 163:19:@16599.4]
  assign storeAddrNotKnownFlags_8_1 = _T_16802 & entriesToCheck_8_1; // @[LoadQueue.scala 163:19:@16601.4]
  assign storeAddrNotKnownFlags_8_2 = _T_16805 & entriesToCheck_8_2; // @[LoadQueue.scala 163:19:@16603.4]
  assign storeAddrNotKnownFlags_8_3 = _T_16808 & entriesToCheck_8_3; // @[LoadQueue.scala 163:19:@16605.4]
  assign storeAddrNotKnownFlags_8_4 = _T_16811 & entriesToCheck_8_4; // @[LoadQueue.scala 163:19:@16607.4]
  assign storeAddrNotKnownFlags_8_5 = _T_16814 & entriesToCheck_8_5; // @[LoadQueue.scala 163:19:@16609.4]
  assign storeAddrNotKnownFlags_8_6 = _T_16817 & entriesToCheck_8_6; // @[LoadQueue.scala 163:19:@16611.4]
  assign storeAddrNotKnownFlags_8_7 = _T_16820 & entriesToCheck_8_7; // @[LoadQueue.scala 163:19:@16613.4]
  assign storeAddrNotKnownFlags_8_8 = _T_16823 & entriesToCheck_8_8; // @[LoadQueue.scala 163:19:@16615.4]
  assign storeAddrNotKnownFlags_8_9 = _T_16826 & entriesToCheck_8_9; // @[LoadQueue.scala 163:19:@16617.4]
  assign storeAddrNotKnownFlags_8_10 = _T_16829 & entriesToCheck_8_10; // @[LoadQueue.scala 163:19:@16619.4]
  assign storeAddrNotKnownFlags_8_11 = _T_16832 & entriesToCheck_8_11; // @[LoadQueue.scala 163:19:@16621.4]
  assign storeAddrNotKnownFlags_8_12 = _T_16835 & entriesToCheck_8_12; // @[LoadQueue.scala 163:19:@16623.4]
  assign storeAddrNotKnownFlags_8_13 = _T_16838 & entriesToCheck_8_13; // @[LoadQueue.scala 163:19:@16625.4]
  assign storeAddrNotKnownFlags_8_14 = _T_16841 & entriesToCheck_8_14; // @[LoadQueue.scala 163:19:@16627.4]
  assign storeAddrNotKnownFlags_8_15 = _T_16844 & entriesToCheck_8_15; // @[LoadQueue.scala 163:19:@16629.4]
  assign storeAddrNotKnownFlags_9_0 = _T_16799 & entriesToCheck_9_0; // @[LoadQueue.scala 163:19:@16647.4]
  assign storeAddrNotKnownFlags_9_1 = _T_16802 & entriesToCheck_9_1; // @[LoadQueue.scala 163:19:@16649.4]
  assign storeAddrNotKnownFlags_9_2 = _T_16805 & entriesToCheck_9_2; // @[LoadQueue.scala 163:19:@16651.4]
  assign storeAddrNotKnownFlags_9_3 = _T_16808 & entriesToCheck_9_3; // @[LoadQueue.scala 163:19:@16653.4]
  assign storeAddrNotKnownFlags_9_4 = _T_16811 & entriesToCheck_9_4; // @[LoadQueue.scala 163:19:@16655.4]
  assign storeAddrNotKnownFlags_9_5 = _T_16814 & entriesToCheck_9_5; // @[LoadQueue.scala 163:19:@16657.4]
  assign storeAddrNotKnownFlags_9_6 = _T_16817 & entriesToCheck_9_6; // @[LoadQueue.scala 163:19:@16659.4]
  assign storeAddrNotKnownFlags_9_7 = _T_16820 & entriesToCheck_9_7; // @[LoadQueue.scala 163:19:@16661.4]
  assign storeAddrNotKnownFlags_9_8 = _T_16823 & entriesToCheck_9_8; // @[LoadQueue.scala 163:19:@16663.4]
  assign storeAddrNotKnownFlags_9_9 = _T_16826 & entriesToCheck_9_9; // @[LoadQueue.scala 163:19:@16665.4]
  assign storeAddrNotKnownFlags_9_10 = _T_16829 & entriesToCheck_9_10; // @[LoadQueue.scala 163:19:@16667.4]
  assign storeAddrNotKnownFlags_9_11 = _T_16832 & entriesToCheck_9_11; // @[LoadQueue.scala 163:19:@16669.4]
  assign storeAddrNotKnownFlags_9_12 = _T_16835 & entriesToCheck_9_12; // @[LoadQueue.scala 163:19:@16671.4]
  assign storeAddrNotKnownFlags_9_13 = _T_16838 & entriesToCheck_9_13; // @[LoadQueue.scala 163:19:@16673.4]
  assign storeAddrNotKnownFlags_9_14 = _T_16841 & entriesToCheck_9_14; // @[LoadQueue.scala 163:19:@16675.4]
  assign storeAddrNotKnownFlags_9_15 = _T_16844 & entriesToCheck_9_15; // @[LoadQueue.scala 163:19:@16677.4]
  assign storeAddrNotKnownFlags_10_0 = _T_16799 & entriesToCheck_10_0; // @[LoadQueue.scala 163:19:@16695.4]
  assign storeAddrNotKnownFlags_10_1 = _T_16802 & entriesToCheck_10_1; // @[LoadQueue.scala 163:19:@16697.4]
  assign storeAddrNotKnownFlags_10_2 = _T_16805 & entriesToCheck_10_2; // @[LoadQueue.scala 163:19:@16699.4]
  assign storeAddrNotKnownFlags_10_3 = _T_16808 & entriesToCheck_10_3; // @[LoadQueue.scala 163:19:@16701.4]
  assign storeAddrNotKnownFlags_10_4 = _T_16811 & entriesToCheck_10_4; // @[LoadQueue.scala 163:19:@16703.4]
  assign storeAddrNotKnownFlags_10_5 = _T_16814 & entriesToCheck_10_5; // @[LoadQueue.scala 163:19:@16705.4]
  assign storeAddrNotKnownFlags_10_6 = _T_16817 & entriesToCheck_10_6; // @[LoadQueue.scala 163:19:@16707.4]
  assign storeAddrNotKnownFlags_10_7 = _T_16820 & entriesToCheck_10_7; // @[LoadQueue.scala 163:19:@16709.4]
  assign storeAddrNotKnownFlags_10_8 = _T_16823 & entriesToCheck_10_8; // @[LoadQueue.scala 163:19:@16711.4]
  assign storeAddrNotKnownFlags_10_9 = _T_16826 & entriesToCheck_10_9; // @[LoadQueue.scala 163:19:@16713.4]
  assign storeAddrNotKnownFlags_10_10 = _T_16829 & entriesToCheck_10_10; // @[LoadQueue.scala 163:19:@16715.4]
  assign storeAddrNotKnownFlags_10_11 = _T_16832 & entriesToCheck_10_11; // @[LoadQueue.scala 163:19:@16717.4]
  assign storeAddrNotKnownFlags_10_12 = _T_16835 & entriesToCheck_10_12; // @[LoadQueue.scala 163:19:@16719.4]
  assign storeAddrNotKnownFlags_10_13 = _T_16838 & entriesToCheck_10_13; // @[LoadQueue.scala 163:19:@16721.4]
  assign storeAddrNotKnownFlags_10_14 = _T_16841 & entriesToCheck_10_14; // @[LoadQueue.scala 163:19:@16723.4]
  assign storeAddrNotKnownFlags_10_15 = _T_16844 & entriesToCheck_10_15; // @[LoadQueue.scala 163:19:@16725.4]
  assign storeAddrNotKnownFlags_11_0 = _T_16799 & entriesToCheck_11_0; // @[LoadQueue.scala 163:19:@16743.4]
  assign storeAddrNotKnownFlags_11_1 = _T_16802 & entriesToCheck_11_1; // @[LoadQueue.scala 163:19:@16745.4]
  assign storeAddrNotKnownFlags_11_2 = _T_16805 & entriesToCheck_11_2; // @[LoadQueue.scala 163:19:@16747.4]
  assign storeAddrNotKnownFlags_11_3 = _T_16808 & entriesToCheck_11_3; // @[LoadQueue.scala 163:19:@16749.4]
  assign storeAddrNotKnownFlags_11_4 = _T_16811 & entriesToCheck_11_4; // @[LoadQueue.scala 163:19:@16751.4]
  assign storeAddrNotKnownFlags_11_5 = _T_16814 & entriesToCheck_11_5; // @[LoadQueue.scala 163:19:@16753.4]
  assign storeAddrNotKnownFlags_11_6 = _T_16817 & entriesToCheck_11_6; // @[LoadQueue.scala 163:19:@16755.4]
  assign storeAddrNotKnownFlags_11_7 = _T_16820 & entriesToCheck_11_7; // @[LoadQueue.scala 163:19:@16757.4]
  assign storeAddrNotKnownFlags_11_8 = _T_16823 & entriesToCheck_11_8; // @[LoadQueue.scala 163:19:@16759.4]
  assign storeAddrNotKnownFlags_11_9 = _T_16826 & entriesToCheck_11_9; // @[LoadQueue.scala 163:19:@16761.4]
  assign storeAddrNotKnownFlags_11_10 = _T_16829 & entriesToCheck_11_10; // @[LoadQueue.scala 163:19:@16763.4]
  assign storeAddrNotKnownFlags_11_11 = _T_16832 & entriesToCheck_11_11; // @[LoadQueue.scala 163:19:@16765.4]
  assign storeAddrNotKnownFlags_11_12 = _T_16835 & entriesToCheck_11_12; // @[LoadQueue.scala 163:19:@16767.4]
  assign storeAddrNotKnownFlags_11_13 = _T_16838 & entriesToCheck_11_13; // @[LoadQueue.scala 163:19:@16769.4]
  assign storeAddrNotKnownFlags_11_14 = _T_16841 & entriesToCheck_11_14; // @[LoadQueue.scala 163:19:@16771.4]
  assign storeAddrNotKnownFlags_11_15 = _T_16844 & entriesToCheck_11_15; // @[LoadQueue.scala 163:19:@16773.4]
  assign storeAddrNotKnownFlags_12_0 = _T_16799 & entriesToCheck_12_0; // @[LoadQueue.scala 163:19:@16791.4]
  assign storeAddrNotKnownFlags_12_1 = _T_16802 & entriesToCheck_12_1; // @[LoadQueue.scala 163:19:@16793.4]
  assign storeAddrNotKnownFlags_12_2 = _T_16805 & entriesToCheck_12_2; // @[LoadQueue.scala 163:19:@16795.4]
  assign storeAddrNotKnownFlags_12_3 = _T_16808 & entriesToCheck_12_3; // @[LoadQueue.scala 163:19:@16797.4]
  assign storeAddrNotKnownFlags_12_4 = _T_16811 & entriesToCheck_12_4; // @[LoadQueue.scala 163:19:@16799.4]
  assign storeAddrNotKnownFlags_12_5 = _T_16814 & entriesToCheck_12_5; // @[LoadQueue.scala 163:19:@16801.4]
  assign storeAddrNotKnownFlags_12_6 = _T_16817 & entriesToCheck_12_6; // @[LoadQueue.scala 163:19:@16803.4]
  assign storeAddrNotKnownFlags_12_7 = _T_16820 & entriesToCheck_12_7; // @[LoadQueue.scala 163:19:@16805.4]
  assign storeAddrNotKnownFlags_12_8 = _T_16823 & entriesToCheck_12_8; // @[LoadQueue.scala 163:19:@16807.4]
  assign storeAddrNotKnownFlags_12_9 = _T_16826 & entriesToCheck_12_9; // @[LoadQueue.scala 163:19:@16809.4]
  assign storeAddrNotKnownFlags_12_10 = _T_16829 & entriesToCheck_12_10; // @[LoadQueue.scala 163:19:@16811.4]
  assign storeAddrNotKnownFlags_12_11 = _T_16832 & entriesToCheck_12_11; // @[LoadQueue.scala 163:19:@16813.4]
  assign storeAddrNotKnownFlags_12_12 = _T_16835 & entriesToCheck_12_12; // @[LoadQueue.scala 163:19:@16815.4]
  assign storeAddrNotKnownFlags_12_13 = _T_16838 & entriesToCheck_12_13; // @[LoadQueue.scala 163:19:@16817.4]
  assign storeAddrNotKnownFlags_12_14 = _T_16841 & entriesToCheck_12_14; // @[LoadQueue.scala 163:19:@16819.4]
  assign storeAddrNotKnownFlags_12_15 = _T_16844 & entriesToCheck_12_15; // @[LoadQueue.scala 163:19:@16821.4]
  assign storeAddrNotKnownFlags_13_0 = _T_16799 & entriesToCheck_13_0; // @[LoadQueue.scala 163:19:@16839.4]
  assign storeAddrNotKnownFlags_13_1 = _T_16802 & entriesToCheck_13_1; // @[LoadQueue.scala 163:19:@16841.4]
  assign storeAddrNotKnownFlags_13_2 = _T_16805 & entriesToCheck_13_2; // @[LoadQueue.scala 163:19:@16843.4]
  assign storeAddrNotKnownFlags_13_3 = _T_16808 & entriesToCheck_13_3; // @[LoadQueue.scala 163:19:@16845.4]
  assign storeAddrNotKnownFlags_13_4 = _T_16811 & entriesToCheck_13_4; // @[LoadQueue.scala 163:19:@16847.4]
  assign storeAddrNotKnownFlags_13_5 = _T_16814 & entriesToCheck_13_5; // @[LoadQueue.scala 163:19:@16849.4]
  assign storeAddrNotKnownFlags_13_6 = _T_16817 & entriesToCheck_13_6; // @[LoadQueue.scala 163:19:@16851.4]
  assign storeAddrNotKnownFlags_13_7 = _T_16820 & entriesToCheck_13_7; // @[LoadQueue.scala 163:19:@16853.4]
  assign storeAddrNotKnownFlags_13_8 = _T_16823 & entriesToCheck_13_8; // @[LoadQueue.scala 163:19:@16855.4]
  assign storeAddrNotKnownFlags_13_9 = _T_16826 & entriesToCheck_13_9; // @[LoadQueue.scala 163:19:@16857.4]
  assign storeAddrNotKnownFlags_13_10 = _T_16829 & entriesToCheck_13_10; // @[LoadQueue.scala 163:19:@16859.4]
  assign storeAddrNotKnownFlags_13_11 = _T_16832 & entriesToCheck_13_11; // @[LoadQueue.scala 163:19:@16861.4]
  assign storeAddrNotKnownFlags_13_12 = _T_16835 & entriesToCheck_13_12; // @[LoadQueue.scala 163:19:@16863.4]
  assign storeAddrNotKnownFlags_13_13 = _T_16838 & entriesToCheck_13_13; // @[LoadQueue.scala 163:19:@16865.4]
  assign storeAddrNotKnownFlags_13_14 = _T_16841 & entriesToCheck_13_14; // @[LoadQueue.scala 163:19:@16867.4]
  assign storeAddrNotKnownFlags_13_15 = _T_16844 & entriesToCheck_13_15; // @[LoadQueue.scala 163:19:@16869.4]
  assign storeAddrNotKnownFlags_14_0 = _T_16799 & entriesToCheck_14_0; // @[LoadQueue.scala 163:19:@16887.4]
  assign storeAddrNotKnownFlags_14_1 = _T_16802 & entriesToCheck_14_1; // @[LoadQueue.scala 163:19:@16889.4]
  assign storeAddrNotKnownFlags_14_2 = _T_16805 & entriesToCheck_14_2; // @[LoadQueue.scala 163:19:@16891.4]
  assign storeAddrNotKnownFlags_14_3 = _T_16808 & entriesToCheck_14_3; // @[LoadQueue.scala 163:19:@16893.4]
  assign storeAddrNotKnownFlags_14_4 = _T_16811 & entriesToCheck_14_4; // @[LoadQueue.scala 163:19:@16895.4]
  assign storeAddrNotKnownFlags_14_5 = _T_16814 & entriesToCheck_14_5; // @[LoadQueue.scala 163:19:@16897.4]
  assign storeAddrNotKnownFlags_14_6 = _T_16817 & entriesToCheck_14_6; // @[LoadQueue.scala 163:19:@16899.4]
  assign storeAddrNotKnownFlags_14_7 = _T_16820 & entriesToCheck_14_7; // @[LoadQueue.scala 163:19:@16901.4]
  assign storeAddrNotKnownFlags_14_8 = _T_16823 & entriesToCheck_14_8; // @[LoadQueue.scala 163:19:@16903.4]
  assign storeAddrNotKnownFlags_14_9 = _T_16826 & entriesToCheck_14_9; // @[LoadQueue.scala 163:19:@16905.4]
  assign storeAddrNotKnownFlags_14_10 = _T_16829 & entriesToCheck_14_10; // @[LoadQueue.scala 163:19:@16907.4]
  assign storeAddrNotKnownFlags_14_11 = _T_16832 & entriesToCheck_14_11; // @[LoadQueue.scala 163:19:@16909.4]
  assign storeAddrNotKnownFlags_14_12 = _T_16835 & entriesToCheck_14_12; // @[LoadQueue.scala 163:19:@16911.4]
  assign storeAddrNotKnownFlags_14_13 = _T_16838 & entriesToCheck_14_13; // @[LoadQueue.scala 163:19:@16913.4]
  assign storeAddrNotKnownFlags_14_14 = _T_16841 & entriesToCheck_14_14; // @[LoadQueue.scala 163:19:@16915.4]
  assign storeAddrNotKnownFlags_14_15 = _T_16844 & entriesToCheck_14_15; // @[LoadQueue.scala 163:19:@16917.4]
  assign storeAddrNotKnownFlags_15_0 = _T_16799 & entriesToCheck_15_0; // @[LoadQueue.scala 163:19:@16935.4]
  assign storeAddrNotKnownFlags_15_1 = _T_16802 & entriesToCheck_15_1; // @[LoadQueue.scala 163:19:@16937.4]
  assign storeAddrNotKnownFlags_15_2 = _T_16805 & entriesToCheck_15_2; // @[LoadQueue.scala 163:19:@16939.4]
  assign storeAddrNotKnownFlags_15_3 = _T_16808 & entriesToCheck_15_3; // @[LoadQueue.scala 163:19:@16941.4]
  assign storeAddrNotKnownFlags_15_4 = _T_16811 & entriesToCheck_15_4; // @[LoadQueue.scala 163:19:@16943.4]
  assign storeAddrNotKnownFlags_15_5 = _T_16814 & entriesToCheck_15_5; // @[LoadQueue.scala 163:19:@16945.4]
  assign storeAddrNotKnownFlags_15_6 = _T_16817 & entriesToCheck_15_6; // @[LoadQueue.scala 163:19:@16947.4]
  assign storeAddrNotKnownFlags_15_7 = _T_16820 & entriesToCheck_15_7; // @[LoadQueue.scala 163:19:@16949.4]
  assign storeAddrNotKnownFlags_15_8 = _T_16823 & entriesToCheck_15_8; // @[LoadQueue.scala 163:19:@16951.4]
  assign storeAddrNotKnownFlags_15_9 = _T_16826 & entriesToCheck_15_9; // @[LoadQueue.scala 163:19:@16953.4]
  assign storeAddrNotKnownFlags_15_10 = _T_16829 & entriesToCheck_15_10; // @[LoadQueue.scala 163:19:@16955.4]
  assign storeAddrNotKnownFlags_15_11 = _T_16832 & entriesToCheck_15_11; // @[LoadQueue.scala 163:19:@16957.4]
  assign storeAddrNotKnownFlags_15_12 = _T_16835 & entriesToCheck_15_12; // @[LoadQueue.scala 163:19:@16959.4]
  assign storeAddrNotKnownFlags_15_13 = _T_16838 & entriesToCheck_15_13; // @[LoadQueue.scala 163:19:@16961.4]
  assign storeAddrNotKnownFlags_15_14 = _T_16841 & entriesToCheck_15_14; // @[LoadQueue.scala 163:19:@16963.4]
  assign storeAddrNotKnownFlags_15_15 = _T_16844 & entriesToCheck_15_15; // @[LoadQueue.scala 163:19:@16965.4]
  assign _T_18002 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@17296.4]
  assign _T_18009 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8}; // @[Mux.scala 19:72:@17303.4]
  assign _T_18010 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,_T_18002}; // @[Mux.scala 19:72:@17304.4]
  assign _T_18012 = _T_2689 ? _T_18010 : 16'h0; // @[Mux.scala 19:72:@17305.4]
  assign _T_18019 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@17312.4]
  assign _T_18026 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9}; // @[Mux.scala 19:72:@17319.4]
  assign _T_18027 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,_T_18019}; // @[Mux.scala 19:72:@17320.4]
  assign _T_18029 = _T_2690 ? _T_18027 : 16'h0; // @[Mux.scala 19:72:@17321.4]
  assign _T_18036 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@17328.4]
  assign _T_18043 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10}; // @[Mux.scala 19:72:@17335.4]
  assign _T_18044 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,_T_18036}; // @[Mux.scala 19:72:@17336.4]
  assign _T_18046 = _T_2691 ? _T_18044 : 16'h0; // @[Mux.scala 19:72:@17337.4]
  assign _T_18053 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@17344.4]
  assign _T_18060 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11}; // @[Mux.scala 19:72:@17351.4]
  assign _T_18061 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,_T_18053}; // @[Mux.scala 19:72:@17352.4]
  assign _T_18063 = _T_2692 ? _T_18061 : 16'h0; // @[Mux.scala 19:72:@17353.4]
  assign _T_18070 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@17360.4]
  assign _T_18077 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12}; // @[Mux.scala 19:72:@17367.4]
  assign _T_18078 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,_T_18070}; // @[Mux.scala 19:72:@17368.4]
  assign _T_18080 = _T_2693 ? _T_18078 : 16'h0; // @[Mux.scala 19:72:@17369.4]
  assign _T_18087 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@17376.4]
  assign _T_18094 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13}; // @[Mux.scala 19:72:@17383.4]
  assign _T_18095 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,_T_18087}; // @[Mux.scala 19:72:@17384.4]
  assign _T_18097 = _T_2694 ? _T_18095 : 16'h0; // @[Mux.scala 19:72:@17385.4]
  assign _T_18104 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@17392.4]
  assign _T_18111 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14}; // @[Mux.scala 19:72:@17399.4]
  assign _T_18112 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,_T_18104}; // @[Mux.scala 19:72:@17400.4]
  assign _T_18114 = _T_2695 ? _T_18112 : 16'h0; // @[Mux.scala 19:72:@17401.4]
  assign _T_18121 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7}; // @[Mux.scala 19:72:@17408.4]
  assign _T_18128 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15}; // @[Mux.scala 19:72:@17415.4]
  assign _T_18129 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,_T_18121}; // @[Mux.scala 19:72:@17416.4]
  assign _T_18131 = _T_2696 ? _T_18129 : 16'h0; // @[Mux.scala 19:72:@17417.4]
  assign _T_18146 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,_T_18009}; // @[Mux.scala 19:72:@17432.4]
  assign _T_18148 = _T_2697 ? _T_18146 : 16'h0; // @[Mux.scala 19:72:@17433.4]
  assign _T_18163 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,_T_18026}; // @[Mux.scala 19:72:@17448.4]
  assign _T_18165 = _T_2698 ? _T_18163 : 16'h0; // @[Mux.scala 19:72:@17449.4]
  assign _T_18180 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,_T_18043}; // @[Mux.scala 19:72:@17464.4]
  assign _T_18182 = _T_2699 ? _T_18180 : 16'h0; // @[Mux.scala 19:72:@17465.4]
  assign _T_18197 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,_T_18060}; // @[Mux.scala 19:72:@17480.4]
  assign _T_18199 = _T_2700 ? _T_18197 : 16'h0; // @[Mux.scala 19:72:@17481.4]
  assign _T_18214 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,_T_18077}; // @[Mux.scala 19:72:@17496.4]
  assign _T_18216 = _T_2701 ? _T_18214 : 16'h0; // @[Mux.scala 19:72:@17497.4]
  assign _T_18231 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,_T_18094}; // @[Mux.scala 19:72:@17512.4]
  assign _T_18233 = _T_2702 ? _T_18231 : 16'h0; // @[Mux.scala 19:72:@17513.4]
  assign _T_18248 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,_T_18111}; // @[Mux.scala 19:72:@17528.4]
  assign _T_18250 = _T_2703 ? _T_18248 : 16'h0; // @[Mux.scala 19:72:@17529.4]
  assign _T_18265 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,_T_18128}; // @[Mux.scala 19:72:@17544.4]
  assign _T_18267 = _T_2704 ? _T_18265 : 16'h0; // @[Mux.scala 19:72:@17545.4]
  assign _T_18268 = _T_18012 | _T_18029; // @[Mux.scala 19:72:@17546.4]
  assign _T_18269 = _T_18268 | _T_18046; // @[Mux.scala 19:72:@17547.4]
  assign _T_18270 = _T_18269 | _T_18063; // @[Mux.scala 19:72:@17548.4]
  assign _T_18271 = _T_18270 | _T_18080; // @[Mux.scala 19:72:@17549.4]
  assign _T_18272 = _T_18271 | _T_18097; // @[Mux.scala 19:72:@17550.4]
  assign _T_18273 = _T_18272 | _T_18114; // @[Mux.scala 19:72:@17551.4]
  assign _T_18274 = _T_18273 | _T_18131; // @[Mux.scala 19:72:@17552.4]
  assign _T_18275 = _T_18274 | _T_18148; // @[Mux.scala 19:72:@17553.4]
  assign _T_18276 = _T_18275 | _T_18165; // @[Mux.scala 19:72:@17554.4]
  assign _T_18277 = _T_18276 | _T_18182; // @[Mux.scala 19:72:@17555.4]
  assign _T_18278 = _T_18277 | _T_18199; // @[Mux.scala 19:72:@17556.4]
  assign _T_18279 = _T_18278 | _T_18216; // @[Mux.scala 19:72:@17557.4]
  assign _T_18280 = _T_18279 | _T_18233; // @[Mux.scala 19:72:@17558.4]
  assign _T_18281 = _T_18280 | _T_18250; // @[Mux.scala 19:72:@17559.4]
  assign _T_18282 = _T_18281 | _T_18267; // @[Mux.scala 19:72:@17560.4]
  assign _T_18860 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@17910.4]
  assign _T_18867 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8}; // @[Mux.scala 19:72:@17917.4]
  assign _T_18868 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,_T_18860}; // @[Mux.scala 19:72:@17918.4]
  assign _T_18870 = _T_2689 ? _T_18868 : 16'h0; // @[Mux.scala 19:72:@17919.4]
  assign _T_18877 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@17926.4]
  assign _T_18884 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9}; // @[Mux.scala 19:72:@17933.4]
  assign _T_18885 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,_T_18877}; // @[Mux.scala 19:72:@17934.4]
  assign _T_18887 = _T_2690 ? _T_18885 : 16'h0; // @[Mux.scala 19:72:@17935.4]
  assign _T_18894 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@17942.4]
  assign _T_18901 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10}; // @[Mux.scala 19:72:@17949.4]
  assign _T_18902 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,_T_18894}; // @[Mux.scala 19:72:@17950.4]
  assign _T_18904 = _T_2691 ? _T_18902 : 16'h0; // @[Mux.scala 19:72:@17951.4]
  assign _T_18911 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@17958.4]
  assign _T_18918 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11}; // @[Mux.scala 19:72:@17965.4]
  assign _T_18919 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,_T_18911}; // @[Mux.scala 19:72:@17966.4]
  assign _T_18921 = _T_2692 ? _T_18919 : 16'h0; // @[Mux.scala 19:72:@17967.4]
  assign _T_18928 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@17974.4]
  assign _T_18935 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12}; // @[Mux.scala 19:72:@17981.4]
  assign _T_18936 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,_T_18928}; // @[Mux.scala 19:72:@17982.4]
  assign _T_18938 = _T_2693 ? _T_18936 : 16'h0; // @[Mux.scala 19:72:@17983.4]
  assign _T_18945 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@17990.4]
  assign _T_18952 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13}; // @[Mux.scala 19:72:@17997.4]
  assign _T_18953 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,_T_18945}; // @[Mux.scala 19:72:@17998.4]
  assign _T_18955 = _T_2694 ? _T_18953 : 16'h0; // @[Mux.scala 19:72:@17999.4]
  assign _T_18962 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@18006.4]
  assign _T_18969 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14}; // @[Mux.scala 19:72:@18013.4]
  assign _T_18970 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,_T_18962}; // @[Mux.scala 19:72:@18014.4]
  assign _T_18972 = _T_2695 ? _T_18970 : 16'h0; // @[Mux.scala 19:72:@18015.4]
  assign _T_18979 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7}; // @[Mux.scala 19:72:@18022.4]
  assign _T_18986 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15}; // @[Mux.scala 19:72:@18029.4]
  assign _T_18987 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,_T_18979}; // @[Mux.scala 19:72:@18030.4]
  assign _T_18989 = _T_2696 ? _T_18987 : 16'h0; // @[Mux.scala 19:72:@18031.4]
  assign _T_19004 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,_T_18867}; // @[Mux.scala 19:72:@18046.4]
  assign _T_19006 = _T_2697 ? _T_19004 : 16'h0; // @[Mux.scala 19:72:@18047.4]
  assign _T_19021 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,_T_18884}; // @[Mux.scala 19:72:@18062.4]
  assign _T_19023 = _T_2698 ? _T_19021 : 16'h0; // @[Mux.scala 19:72:@18063.4]
  assign _T_19038 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,_T_18901}; // @[Mux.scala 19:72:@18078.4]
  assign _T_19040 = _T_2699 ? _T_19038 : 16'h0; // @[Mux.scala 19:72:@18079.4]
  assign _T_19055 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,_T_18918}; // @[Mux.scala 19:72:@18094.4]
  assign _T_19057 = _T_2700 ? _T_19055 : 16'h0; // @[Mux.scala 19:72:@18095.4]
  assign _T_19072 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,_T_18935}; // @[Mux.scala 19:72:@18110.4]
  assign _T_19074 = _T_2701 ? _T_19072 : 16'h0; // @[Mux.scala 19:72:@18111.4]
  assign _T_19089 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,_T_18952}; // @[Mux.scala 19:72:@18126.4]
  assign _T_19091 = _T_2702 ? _T_19089 : 16'h0; // @[Mux.scala 19:72:@18127.4]
  assign _T_19106 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,_T_18969}; // @[Mux.scala 19:72:@18142.4]
  assign _T_19108 = _T_2703 ? _T_19106 : 16'h0; // @[Mux.scala 19:72:@18143.4]
  assign _T_19123 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,_T_18986}; // @[Mux.scala 19:72:@18158.4]
  assign _T_19125 = _T_2704 ? _T_19123 : 16'h0; // @[Mux.scala 19:72:@18159.4]
  assign _T_19126 = _T_18870 | _T_18887; // @[Mux.scala 19:72:@18160.4]
  assign _T_19127 = _T_19126 | _T_18904; // @[Mux.scala 19:72:@18161.4]
  assign _T_19128 = _T_19127 | _T_18921; // @[Mux.scala 19:72:@18162.4]
  assign _T_19129 = _T_19128 | _T_18938; // @[Mux.scala 19:72:@18163.4]
  assign _T_19130 = _T_19129 | _T_18955; // @[Mux.scala 19:72:@18164.4]
  assign _T_19131 = _T_19130 | _T_18972; // @[Mux.scala 19:72:@18165.4]
  assign _T_19132 = _T_19131 | _T_18989; // @[Mux.scala 19:72:@18166.4]
  assign _T_19133 = _T_19132 | _T_19006; // @[Mux.scala 19:72:@18167.4]
  assign _T_19134 = _T_19133 | _T_19023; // @[Mux.scala 19:72:@18168.4]
  assign _T_19135 = _T_19134 | _T_19040; // @[Mux.scala 19:72:@18169.4]
  assign _T_19136 = _T_19135 | _T_19057; // @[Mux.scala 19:72:@18170.4]
  assign _T_19137 = _T_19136 | _T_19074; // @[Mux.scala 19:72:@18171.4]
  assign _T_19138 = _T_19137 | _T_19091; // @[Mux.scala 19:72:@18172.4]
  assign _T_19139 = _T_19138 | _T_19108; // @[Mux.scala 19:72:@18173.4]
  assign _T_19140 = _T_19139 | _T_19125; // @[Mux.scala 19:72:@18174.4]
  assign _T_19718 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@18524.4]
  assign _T_19725 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8}; // @[Mux.scala 19:72:@18531.4]
  assign _T_19726 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,_T_19718}; // @[Mux.scala 19:72:@18532.4]
  assign _T_19728 = _T_2689 ? _T_19726 : 16'h0; // @[Mux.scala 19:72:@18533.4]
  assign _T_19735 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@18540.4]
  assign _T_19742 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9}; // @[Mux.scala 19:72:@18547.4]
  assign _T_19743 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,_T_19735}; // @[Mux.scala 19:72:@18548.4]
  assign _T_19745 = _T_2690 ? _T_19743 : 16'h0; // @[Mux.scala 19:72:@18549.4]
  assign _T_19752 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@18556.4]
  assign _T_19759 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10}; // @[Mux.scala 19:72:@18563.4]
  assign _T_19760 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,_T_19752}; // @[Mux.scala 19:72:@18564.4]
  assign _T_19762 = _T_2691 ? _T_19760 : 16'h0; // @[Mux.scala 19:72:@18565.4]
  assign _T_19769 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@18572.4]
  assign _T_19776 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11}; // @[Mux.scala 19:72:@18579.4]
  assign _T_19777 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,_T_19769}; // @[Mux.scala 19:72:@18580.4]
  assign _T_19779 = _T_2692 ? _T_19777 : 16'h0; // @[Mux.scala 19:72:@18581.4]
  assign _T_19786 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@18588.4]
  assign _T_19793 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12}; // @[Mux.scala 19:72:@18595.4]
  assign _T_19794 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,_T_19786}; // @[Mux.scala 19:72:@18596.4]
  assign _T_19796 = _T_2693 ? _T_19794 : 16'h0; // @[Mux.scala 19:72:@18597.4]
  assign _T_19803 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@18604.4]
  assign _T_19810 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13}; // @[Mux.scala 19:72:@18611.4]
  assign _T_19811 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,_T_19803}; // @[Mux.scala 19:72:@18612.4]
  assign _T_19813 = _T_2694 ? _T_19811 : 16'h0; // @[Mux.scala 19:72:@18613.4]
  assign _T_19820 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@18620.4]
  assign _T_19827 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14}; // @[Mux.scala 19:72:@18627.4]
  assign _T_19828 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,_T_19820}; // @[Mux.scala 19:72:@18628.4]
  assign _T_19830 = _T_2695 ? _T_19828 : 16'h0; // @[Mux.scala 19:72:@18629.4]
  assign _T_19837 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7}; // @[Mux.scala 19:72:@18636.4]
  assign _T_19844 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15}; // @[Mux.scala 19:72:@18643.4]
  assign _T_19845 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,_T_19837}; // @[Mux.scala 19:72:@18644.4]
  assign _T_19847 = _T_2696 ? _T_19845 : 16'h0; // @[Mux.scala 19:72:@18645.4]
  assign _T_19862 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,_T_19725}; // @[Mux.scala 19:72:@18660.4]
  assign _T_19864 = _T_2697 ? _T_19862 : 16'h0; // @[Mux.scala 19:72:@18661.4]
  assign _T_19879 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,_T_19742}; // @[Mux.scala 19:72:@18676.4]
  assign _T_19881 = _T_2698 ? _T_19879 : 16'h0; // @[Mux.scala 19:72:@18677.4]
  assign _T_19896 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,_T_19759}; // @[Mux.scala 19:72:@18692.4]
  assign _T_19898 = _T_2699 ? _T_19896 : 16'h0; // @[Mux.scala 19:72:@18693.4]
  assign _T_19913 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,_T_19776}; // @[Mux.scala 19:72:@18708.4]
  assign _T_19915 = _T_2700 ? _T_19913 : 16'h0; // @[Mux.scala 19:72:@18709.4]
  assign _T_19930 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,_T_19793}; // @[Mux.scala 19:72:@18724.4]
  assign _T_19932 = _T_2701 ? _T_19930 : 16'h0; // @[Mux.scala 19:72:@18725.4]
  assign _T_19947 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,_T_19810}; // @[Mux.scala 19:72:@18740.4]
  assign _T_19949 = _T_2702 ? _T_19947 : 16'h0; // @[Mux.scala 19:72:@18741.4]
  assign _T_19964 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,_T_19827}; // @[Mux.scala 19:72:@18756.4]
  assign _T_19966 = _T_2703 ? _T_19964 : 16'h0; // @[Mux.scala 19:72:@18757.4]
  assign _T_19981 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,_T_19844}; // @[Mux.scala 19:72:@18772.4]
  assign _T_19983 = _T_2704 ? _T_19981 : 16'h0; // @[Mux.scala 19:72:@18773.4]
  assign _T_19984 = _T_19728 | _T_19745; // @[Mux.scala 19:72:@18774.4]
  assign _T_19985 = _T_19984 | _T_19762; // @[Mux.scala 19:72:@18775.4]
  assign _T_19986 = _T_19985 | _T_19779; // @[Mux.scala 19:72:@18776.4]
  assign _T_19987 = _T_19986 | _T_19796; // @[Mux.scala 19:72:@18777.4]
  assign _T_19988 = _T_19987 | _T_19813; // @[Mux.scala 19:72:@18778.4]
  assign _T_19989 = _T_19988 | _T_19830; // @[Mux.scala 19:72:@18779.4]
  assign _T_19990 = _T_19989 | _T_19847; // @[Mux.scala 19:72:@18780.4]
  assign _T_19991 = _T_19990 | _T_19864; // @[Mux.scala 19:72:@18781.4]
  assign _T_19992 = _T_19991 | _T_19881; // @[Mux.scala 19:72:@18782.4]
  assign _T_19993 = _T_19992 | _T_19898; // @[Mux.scala 19:72:@18783.4]
  assign _T_19994 = _T_19993 | _T_19915; // @[Mux.scala 19:72:@18784.4]
  assign _T_19995 = _T_19994 | _T_19932; // @[Mux.scala 19:72:@18785.4]
  assign _T_19996 = _T_19995 | _T_19949; // @[Mux.scala 19:72:@18786.4]
  assign _T_19997 = _T_19996 | _T_19966; // @[Mux.scala 19:72:@18787.4]
  assign _T_19998 = _T_19997 | _T_19983; // @[Mux.scala 19:72:@18788.4]
  assign _T_20576 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@19138.4]
  assign _T_20583 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8}; // @[Mux.scala 19:72:@19145.4]
  assign _T_20584 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,_T_20576}; // @[Mux.scala 19:72:@19146.4]
  assign _T_20586 = _T_2689 ? _T_20584 : 16'h0; // @[Mux.scala 19:72:@19147.4]
  assign _T_20593 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@19154.4]
  assign _T_20600 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9}; // @[Mux.scala 19:72:@19161.4]
  assign _T_20601 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,_T_20593}; // @[Mux.scala 19:72:@19162.4]
  assign _T_20603 = _T_2690 ? _T_20601 : 16'h0; // @[Mux.scala 19:72:@19163.4]
  assign _T_20610 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@19170.4]
  assign _T_20617 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10}; // @[Mux.scala 19:72:@19177.4]
  assign _T_20618 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,_T_20610}; // @[Mux.scala 19:72:@19178.4]
  assign _T_20620 = _T_2691 ? _T_20618 : 16'h0; // @[Mux.scala 19:72:@19179.4]
  assign _T_20627 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@19186.4]
  assign _T_20634 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11}; // @[Mux.scala 19:72:@19193.4]
  assign _T_20635 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,_T_20627}; // @[Mux.scala 19:72:@19194.4]
  assign _T_20637 = _T_2692 ? _T_20635 : 16'h0; // @[Mux.scala 19:72:@19195.4]
  assign _T_20644 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@19202.4]
  assign _T_20651 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12}; // @[Mux.scala 19:72:@19209.4]
  assign _T_20652 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,_T_20644}; // @[Mux.scala 19:72:@19210.4]
  assign _T_20654 = _T_2693 ? _T_20652 : 16'h0; // @[Mux.scala 19:72:@19211.4]
  assign _T_20661 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@19218.4]
  assign _T_20668 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13}; // @[Mux.scala 19:72:@19225.4]
  assign _T_20669 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,_T_20661}; // @[Mux.scala 19:72:@19226.4]
  assign _T_20671 = _T_2694 ? _T_20669 : 16'h0; // @[Mux.scala 19:72:@19227.4]
  assign _T_20678 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@19234.4]
  assign _T_20685 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14}; // @[Mux.scala 19:72:@19241.4]
  assign _T_20686 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,_T_20678}; // @[Mux.scala 19:72:@19242.4]
  assign _T_20688 = _T_2695 ? _T_20686 : 16'h0; // @[Mux.scala 19:72:@19243.4]
  assign _T_20695 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7}; // @[Mux.scala 19:72:@19250.4]
  assign _T_20702 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15}; // @[Mux.scala 19:72:@19257.4]
  assign _T_20703 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,_T_20695}; // @[Mux.scala 19:72:@19258.4]
  assign _T_20705 = _T_2696 ? _T_20703 : 16'h0; // @[Mux.scala 19:72:@19259.4]
  assign _T_20720 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,_T_20583}; // @[Mux.scala 19:72:@19274.4]
  assign _T_20722 = _T_2697 ? _T_20720 : 16'h0; // @[Mux.scala 19:72:@19275.4]
  assign _T_20737 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,_T_20600}; // @[Mux.scala 19:72:@19290.4]
  assign _T_20739 = _T_2698 ? _T_20737 : 16'h0; // @[Mux.scala 19:72:@19291.4]
  assign _T_20754 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,_T_20617}; // @[Mux.scala 19:72:@19306.4]
  assign _T_20756 = _T_2699 ? _T_20754 : 16'h0; // @[Mux.scala 19:72:@19307.4]
  assign _T_20771 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,_T_20634}; // @[Mux.scala 19:72:@19322.4]
  assign _T_20773 = _T_2700 ? _T_20771 : 16'h0; // @[Mux.scala 19:72:@19323.4]
  assign _T_20788 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,_T_20651}; // @[Mux.scala 19:72:@19338.4]
  assign _T_20790 = _T_2701 ? _T_20788 : 16'h0; // @[Mux.scala 19:72:@19339.4]
  assign _T_20805 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,_T_20668}; // @[Mux.scala 19:72:@19354.4]
  assign _T_20807 = _T_2702 ? _T_20805 : 16'h0; // @[Mux.scala 19:72:@19355.4]
  assign _T_20822 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,_T_20685}; // @[Mux.scala 19:72:@19370.4]
  assign _T_20824 = _T_2703 ? _T_20822 : 16'h0; // @[Mux.scala 19:72:@19371.4]
  assign _T_20839 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,_T_20702}; // @[Mux.scala 19:72:@19386.4]
  assign _T_20841 = _T_2704 ? _T_20839 : 16'h0; // @[Mux.scala 19:72:@19387.4]
  assign _T_20842 = _T_20586 | _T_20603; // @[Mux.scala 19:72:@19388.4]
  assign _T_20843 = _T_20842 | _T_20620; // @[Mux.scala 19:72:@19389.4]
  assign _T_20844 = _T_20843 | _T_20637; // @[Mux.scala 19:72:@19390.4]
  assign _T_20845 = _T_20844 | _T_20654; // @[Mux.scala 19:72:@19391.4]
  assign _T_20846 = _T_20845 | _T_20671; // @[Mux.scala 19:72:@19392.4]
  assign _T_20847 = _T_20846 | _T_20688; // @[Mux.scala 19:72:@19393.4]
  assign _T_20848 = _T_20847 | _T_20705; // @[Mux.scala 19:72:@19394.4]
  assign _T_20849 = _T_20848 | _T_20722; // @[Mux.scala 19:72:@19395.4]
  assign _T_20850 = _T_20849 | _T_20739; // @[Mux.scala 19:72:@19396.4]
  assign _T_20851 = _T_20850 | _T_20756; // @[Mux.scala 19:72:@19397.4]
  assign _T_20852 = _T_20851 | _T_20773; // @[Mux.scala 19:72:@19398.4]
  assign _T_20853 = _T_20852 | _T_20790; // @[Mux.scala 19:72:@19399.4]
  assign _T_20854 = _T_20853 | _T_20807; // @[Mux.scala 19:72:@19400.4]
  assign _T_20855 = _T_20854 | _T_20824; // @[Mux.scala 19:72:@19401.4]
  assign _T_20856 = _T_20855 | _T_20841; // @[Mux.scala 19:72:@19402.4]
  assign _T_21434 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@19752.4]
  assign _T_21441 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8}; // @[Mux.scala 19:72:@19759.4]
  assign _T_21442 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,_T_21434}; // @[Mux.scala 19:72:@19760.4]
  assign _T_21444 = _T_2689 ? _T_21442 : 16'h0; // @[Mux.scala 19:72:@19761.4]
  assign _T_21451 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@19768.4]
  assign _T_21458 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9}; // @[Mux.scala 19:72:@19775.4]
  assign _T_21459 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,_T_21451}; // @[Mux.scala 19:72:@19776.4]
  assign _T_21461 = _T_2690 ? _T_21459 : 16'h0; // @[Mux.scala 19:72:@19777.4]
  assign _T_21468 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@19784.4]
  assign _T_21475 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10}; // @[Mux.scala 19:72:@19791.4]
  assign _T_21476 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,_T_21468}; // @[Mux.scala 19:72:@19792.4]
  assign _T_21478 = _T_2691 ? _T_21476 : 16'h0; // @[Mux.scala 19:72:@19793.4]
  assign _T_21485 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@19800.4]
  assign _T_21492 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11}; // @[Mux.scala 19:72:@19807.4]
  assign _T_21493 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,_T_21485}; // @[Mux.scala 19:72:@19808.4]
  assign _T_21495 = _T_2692 ? _T_21493 : 16'h0; // @[Mux.scala 19:72:@19809.4]
  assign _T_21502 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@19816.4]
  assign _T_21509 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12}; // @[Mux.scala 19:72:@19823.4]
  assign _T_21510 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,_T_21502}; // @[Mux.scala 19:72:@19824.4]
  assign _T_21512 = _T_2693 ? _T_21510 : 16'h0; // @[Mux.scala 19:72:@19825.4]
  assign _T_21519 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@19832.4]
  assign _T_21526 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13}; // @[Mux.scala 19:72:@19839.4]
  assign _T_21527 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,_T_21519}; // @[Mux.scala 19:72:@19840.4]
  assign _T_21529 = _T_2694 ? _T_21527 : 16'h0; // @[Mux.scala 19:72:@19841.4]
  assign _T_21536 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@19848.4]
  assign _T_21543 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14}; // @[Mux.scala 19:72:@19855.4]
  assign _T_21544 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,_T_21536}; // @[Mux.scala 19:72:@19856.4]
  assign _T_21546 = _T_2695 ? _T_21544 : 16'h0; // @[Mux.scala 19:72:@19857.4]
  assign _T_21553 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7}; // @[Mux.scala 19:72:@19864.4]
  assign _T_21560 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15}; // @[Mux.scala 19:72:@19871.4]
  assign _T_21561 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,_T_21553}; // @[Mux.scala 19:72:@19872.4]
  assign _T_21563 = _T_2696 ? _T_21561 : 16'h0; // @[Mux.scala 19:72:@19873.4]
  assign _T_21578 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,_T_21441}; // @[Mux.scala 19:72:@19888.4]
  assign _T_21580 = _T_2697 ? _T_21578 : 16'h0; // @[Mux.scala 19:72:@19889.4]
  assign _T_21595 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,_T_21458}; // @[Mux.scala 19:72:@19904.4]
  assign _T_21597 = _T_2698 ? _T_21595 : 16'h0; // @[Mux.scala 19:72:@19905.4]
  assign _T_21612 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,_T_21475}; // @[Mux.scala 19:72:@19920.4]
  assign _T_21614 = _T_2699 ? _T_21612 : 16'h0; // @[Mux.scala 19:72:@19921.4]
  assign _T_21629 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,_T_21492}; // @[Mux.scala 19:72:@19936.4]
  assign _T_21631 = _T_2700 ? _T_21629 : 16'h0; // @[Mux.scala 19:72:@19937.4]
  assign _T_21646 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,_T_21509}; // @[Mux.scala 19:72:@19952.4]
  assign _T_21648 = _T_2701 ? _T_21646 : 16'h0; // @[Mux.scala 19:72:@19953.4]
  assign _T_21663 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,_T_21526}; // @[Mux.scala 19:72:@19968.4]
  assign _T_21665 = _T_2702 ? _T_21663 : 16'h0; // @[Mux.scala 19:72:@19969.4]
  assign _T_21680 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,_T_21543}; // @[Mux.scala 19:72:@19984.4]
  assign _T_21682 = _T_2703 ? _T_21680 : 16'h0; // @[Mux.scala 19:72:@19985.4]
  assign _T_21697 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,_T_21560}; // @[Mux.scala 19:72:@20000.4]
  assign _T_21699 = _T_2704 ? _T_21697 : 16'h0; // @[Mux.scala 19:72:@20001.4]
  assign _T_21700 = _T_21444 | _T_21461; // @[Mux.scala 19:72:@20002.4]
  assign _T_21701 = _T_21700 | _T_21478; // @[Mux.scala 19:72:@20003.4]
  assign _T_21702 = _T_21701 | _T_21495; // @[Mux.scala 19:72:@20004.4]
  assign _T_21703 = _T_21702 | _T_21512; // @[Mux.scala 19:72:@20005.4]
  assign _T_21704 = _T_21703 | _T_21529; // @[Mux.scala 19:72:@20006.4]
  assign _T_21705 = _T_21704 | _T_21546; // @[Mux.scala 19:72:@20007.4]
  assign _T_21706 = _T_21705 | _T_21563; // @[Mux.scala 19:72:@20008.4]
  assign _T_21707 = _T_21706 | _T_21580; // @[Mux.scala 19:72:@20009.4]
  assign _T_21708 = _T_21707 | _T_21597; // @[Mux.scala 19:72:@20010.4]
  assign _T_21709 = _T_21708 | _T_21614; // @[Mux.scala 19:72:@20011.4]
  assign _T_21710 = _T_21709 | _T_21631; // @[Mux.scala 19:72:@20012.4]
  assign _T_21711 = _T_21710 | _T_21648; // @[Mux.scala 19:72:@20013.4]
  assign _T_21712 = _T_21711 | _T_21665; // @[Mux.scala 19:72:@20014.4]
  assign _T_21713 = _T_21712 | _T_21682; // @[Mux.scala 19:72:@20015.4]
  assign _T_21714 = _T_21713 | _T_21699; // @[Mux.scala 19:72:@20016.4]
  assign _T_22292 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@20366.4]
  assign _T_22299 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8}; // @[Mux.scala 19:72:@20373.4]
  assign _T_22300 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,_T_22292}; // @[Mux.scala 19:72:@20374.4]
  assign _T_22302 = _T_2689 ? _T_22300 : 16'h0; // @[Mux.scala 19:72:@20375.4]
  assign _T_22309 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@20382.4]
  assign _T_22316 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9}; // @[Mux.scala 19:72:@20389.4]
  assign _T_22317 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,_T_22309}; // @[Mux.scala 19:72:@20390.4]
  assign _T_22319 = _T_2690 ? _T_22317 : 16'h0; // @[Mux.scala 19:72:@20391.4]
  assign _T_22326 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@20398.4]
  assign _T_22333 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10}; // @[Mux.scala 19:72:@20405.4]
  assign _T_22334 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,_T_22326}; // @[Mux.scala 19:72:@20406.4]
  assign _T_22336 = _T_2691 ? _T_22334 : 16'h0; // @[Mux.scala 19:72:@20407.4]
  assign _T_22343 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@20414.4]
  assign _T_22350 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11}; // @[Mux.scala 19:72:@20421.4]
  assign _T_22351 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,_T_22343}; // @[Mux.scala 19:72:@20422.4]
  assign _T_22353 = _T_2692 ? _T_22351 : 16'h0; // @[Mux.scala 19:72:@20423.4]
  assign _T_22360 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@20430.4]
  assign _T_22367 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12}; // @[Mux.scala 19:72:@20437.4]
  assign _T_22368 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,_T_22360}; // @[Mux.scala 19:72:@20438.4]
  assign _T_22370 = _T_2693 ? _T_22368 : 16'h0; // @[Mux.scala 19:72:@20439.4]
  assign _T_22377 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@20446.4]
  assign _T_22384 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13}; // @[Mux.scala 19:72:@20453.4]
  assign _T_22385 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,_T_22377}; // @[Mux.scala 19:72:@20454.4]
  assign _T_22387 = _T_2694 ? _T_22385 : 16'h0; // @[Mux.scala 19:72:@20455.4]
  assign _T_22394 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@20462.4]
  assign _T_22401 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14}; // @[Mux.scala 19:72:@20469.4]
  assign _T_22402 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,_T_22394}; // @[Mux.scala 19:72:@20470.4]
  assign _T_22404 = _T_2695 ? _T_22402 : 16'h0; // @[Mux.scala 19:72:@20471.4]
  assign _T_22411 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7}; // @[Mux.scala 19:72:@20478.4]
  assign _T_22418 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15}; // @[Mux.scala 19:72:@20485.4]
  assign _T_22419 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,_T_22411}; // @[Mux.scala 19:72:@20486.4]
  assign _T_22421 = _T_2696 ? _T_22419 : 16'h0; // @[Mux.scala 19:72:@20487.4]
  assign _T_22436 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,_T_22299}; // @[Mux.scala 19:72:@20502.4]
  assign _T_22438 = _T_2697 ? _T_22436 : 16'h0; // @[Mux.scala 19:72:@20503.4]
  assign _T_22453 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,_T_22316}; // @[Mux.scala 19:72:@20518.4]
  assign _T_22455 = _T_2698 ? _T_22453 : 16'h0; // @[Mux.scala 19:72:@20519.4]
  assign _T_22470 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,_T_22333}; // @[Mux.scala 19:72:@20534.4]
  assign _T_22472 = _T_2699 ? _T_22470 : 16'h0; // @[Mux.scala 19:72:@20535.4]
  assign _T_22487 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,_T_22350}; // @[Mux.scala 19:72:@20550.4]
  assign _T_22489 = _T_2700 ? _T_22487 : 16'h0; // @[Mux.scala 19:72:@20551.4]
  assign _T_22504 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,_T_22367}; // @[Mux.scala 19:72:@20566.4]
  assign _T_22506 = _T_2701 ? _T_22504 : 16'h0; // @[Mux.scala 19:72:@20567.4]
  assign _T_22521 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,_T_22384}; // @[Mux.scala 19:72:@20582.4]
  assign _T_22523 = _T_2702 ? _T_22521 : 16'h0; // @[Mux.scala 19:72:@20583.4]
  assign _T_22538 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,_T_22401}; // @[Mux.scala 19:72:@20598.4]
  assign _T_22540 = _T_2703 ? _T_22538 : 16'h0; // @[Mux.scala 19:72:@20599.4]
  assign _T_22555 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,_T_22418}; // @[Mux.scala 19:72:@20614.4]
  assign _T_22557 = _T_2704 ? _T_22555 : 16'h0; // @[Mux.scala 19:72:@20615.4]
  assign _T_22558 = _T_22302 | _T_22319; // @[Mux.scala 19:72:@20616.4]
  assign _T_22559 = _T_22558 | _T_22336; // @[Mux.scala 19:72:@20617.4]
  assign _T_22560 = _T_22559 | _T_22353; // @[Mux.scala 19:72:@20618.4]
  assign _T_22561 = _T_22560 | _T_22370; // @[Mux.scala 19:72:@20619.4]
  assign _T_22562 = _T_22561 | _T_22387; // @[Mux.scala 19:72:@20620.4]
  assign _T_22563 = _T_22562 | _T_22404; // @[Mux.scala 19:72:@20621.4]
  assign _T_22564 = _T_22563 | _T_22421; // @[Mux.scala 19:72:@20622.4]
  assign _T_22565 = _T_22564 | _T_22438; // @[Mux.scala 19:72:@20623.4]
  assign _T_22566 = _T_22565 | _T_22455; // @[Mux.scala 19:72:@20624.4]
  assign _T_22567 = _T_22566 | _T_22472; // @[Mux.scala 19:72:@20625.4]
  assign _T_22568 = _T_22567 | _T_22489; // @[Mux.scala 19:72:@20626.4]
  assign _T_22569 = _T_22568 | _T_22506; // @[Mux.scala 19:72:@20627.4]
  assign _T_22570 = _T_22569 | _T_22523; // @[Mux.scala 19:72:@20628.4]
  assign _T_22571 = _T_22570 | _T_22540; // @[Mux.scala 19:72:@20629.4]
  assign _T_22572 = _T_22571 | _T_22557; // @[Mux.scala 19:72:@20630.4]
  assign _T_23150 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@20980.4]
  assign _T_23157 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8}; // @[Mux.scala 19:72:@20987.4]
  assign _T_23158 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,_T_23150}; // @[Mux.scala 19:72:@20988.4]
  assign _T_23160 = _T_2689 ? _T_23158 : 16'h0; // @[Mux.scala 19:72:@20989.4]
  assign _T_23167 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@20996.4]
  assign _T_23174 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9}; // @[Mux.scala 19:72:@21003.4]
  assign _T_23175 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,_T_23167}; // @[Mux.scala 19:72:@21004.4]
  assign _T_23177 = _T_2690 ? _T_23175 : 16'h0; // @[Mux.scala 19:72:@21005.4]
  assign _T_23184 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@21012.4]
  assign _T_23191 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10}; // @[Mux.scala 19:72:@21019.4]
  assign _T_23192 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,_T_23184}; // @[Mux.scala 19:72:@21020.4]
  assign _T_23194 = _T_2691 ? _T_23192 : 16'h0; // @[Mux.scala 19:72:@21021.4]
  assign _T_23201 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@21028.4]
  assign _T_23208 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11}; // @[Mux.scala 19:72:@21035.4]
  assign _T_23209 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,_T_23201}; // @[Mux.scala 19:72:@21036.4]
  assign _T_23211 = _T_2692 ? _T_23209 : 16'h0; // @[Mux.scala 19:72:@21037.4]
  assign _T_23218 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@21044.4]
  assign _T_23225 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12}; // @[Mux.scala 19:72:@21051.4]
  assign _T_23226 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,_T_23218}; // @[Mux.scala 19:72:@21052.4]
  assign _T_23228 = _T_2693 ? _T_23226 : 16'h0; // @[Mux.scala 19:72:@21053.4]
  assign _T_23235 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@21060.4]
  assign _T_23242 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13}; // @[Mux.scala 19:72:@21067.4]
  assign _T_23243 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,_T_23235}; // @[Mux.scala 19:72:@21068.4]
  assign _T_23245 = _T_2694 ? _T_23243 : 16'h0; // @[Mux.scala 19:72:@21069.4]
  assign _T_23252 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@21076.4]
  assign _T_23259 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14}; // @[Mux.scala 19:72:@21083.4]
  assign _T_23260 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,_T_23252}; // @[Mux.scala 19:72:@21084.4]
  assign _T_23262 = _T_2695 ? _T_23260 : 16'h0; // @[Mux.scala 19:72:@21085.4]
  assign _T_23269 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7}; // @[Mux.scala 19:72:@21092.4]
  assign _T_23276 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15}; // @[Mux.scala 19:72:@21099.4]
  assign _T_23277 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,_T_23269}; // @[Mux.scala 19:72:@21100.4]
  assign _T_23279 = _T_2696 ? _T_23277 : 16'h0; // @[Mux.scala 19:72:@21101.4]
  assign _T_23294 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,_T_23157}; // @[Mux.scala 19:72:@21116.4]
  assign _T_23296 = _T_2697 ? _T_23294 : 16'h0; // @[Mux.scala 19:72:@21117.4]
  assign _T_23311 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,_T_23174}; // @[Mux.scala 19:72:@21132.4]
  assign _T_23313 = _T_2698 ? _T_23311 : 16'h0; // @[Mux.scala 19:72:@21133.4]
  assign _T_23328 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,_T_23191}; // @[Mux.scala 19:72:@21148.4]
  assign _T_23330 = _T_2699 ? _T_23328 : 16'h0; // @[Mux.scala 19:72:@21149.4]
  assign _T_23345 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,_T_23208}; // @[Mux.scala 19:72:@21164.4]
  assign _T_23347 = _T_2700 ? _T_23345 : 16'h0; // @[Mux.scala 19:72:@21165.4]
  assign _T_23362 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,_T_23225}; // @[Mux.scala 19:72:@21180.4]
  assign _T_23364 = _T_2701 ? _T_23362 : 16'h0; // @[Mux.scala 19:72:@21181.4]
  assign _T_23379 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,_T_23242}; // @[Mux.scala 19:72:@21196.4]
  assign _T_23381 = _T_2702 ? _T_23379 : 16'h0; // @[Mux.scala 19:72:@21197.4]
  assign _T_23396 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,_T_23259}; // @[Mux.scala 19:72:@21212.4]
  assign _T_23398 = _T_2703 ? _T_23396 : 16'h0; // @[Mux.scala 19:72:@21213.4]
  assign _T_23413 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,_T_23276}; // @[Mux.scala 19:72:@21228.4]
  assign _T_23415 = _T_2704 ? _T_23413 : 16'h0; // @[Mux.scala 19:72:@21229.4]
  assign _T_23416 = _T_23160 | _T_23177; // @[Mux.scala 19:72:@21230.4]
  assign _T_23417 = _T_23416 | _T_23194; // @[Mux.scala 19:72:@21231.4]
  assign _T_23418 = _T_23417 | _T_23211; // @[Mux.scala 19:72:@21232.4]
  assign _T_23419 = _T_23418 | _T_23228; // @[Mux.scala 19:72:@21233.4]
  assign _T_23420 = _T_23419 | _T_23245; // @[Mux.scala 19:72:@21234.4]
  assign _T_23421 = _T_23420 | _T_23262; // @[Mux.scala 19:72:@21235.4]
  assign _T_23422 = _T_23421 | _T_23279; // @[Mux.scala 19:72:@21236.4]
  assign _T_23423 = _T_23422 | _T_23296; // @[Mux.scala 19:72:@21237.4]
  assign _T_23424 = _T_23423 | _T_23313; // @[Mux.scala 19:72:@21238.4]
  assign _T_23425 = _T_23424 | _T_23330; // @[Mux.scala 19:72:@21239.4]
  assign _T_23426 = _T_23425 | _T_23347; // @[Mux.scala 19:72:@21240.4]
  assign _T_23427 = _T_23426 | _T_23364; // @[Mux.scala 19:72:@21241.4]
  assign _T_23428 = _T_23427 | _T_23381; // @[Mux.scala 19:72:@21242.4]
  assign _T_23429 = _T_23428 | _T_23398; // @[Mux.scala 19:72:@21243.4]
  assign _T_23430 = _T_23429 | _T_23415; // @[Mux.scala 19:72:@21244.4]
  assign _T_24008 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@21594.4]
  assign _T_24015 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8}; // @[Mux.scala 19:72:@21601.4]
  assign _T_24016 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,_T_24008}; // @[Mux.scala 19:72:@21602.4]
  assign _T_24018 = _T_2689 ? _T_24016 : 16'h0; // @[Mux.scala 19:72:@21603.4]
  assign _T_24025 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@21610.4]
  assign _T_24032 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9}; // @[Mux.scala 19:72:@21617.4]
  assign _T_24033 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,_T_24025}; // @[Mux.scala 19:72:@21618.4]
  assign _T_24035 = _T_2690 ? _T_24033 : 16'h0; // @[Mux.scala 19:72:@21619.4]
  assign _T_24042 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@21626.4]
  assign _T_24049 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10}; // @[Mux.scala 19:72:@21633.4]
  assign _T_24050 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,_T_24042}; // @[Mux.scala 19:72:@21634.4]
  assign _T_24052 = _T_2691 ? _T_24050 : 16'h0; // @[Mux.scala 19:72:@21635.4]
  assign _T_24059 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@21642.4]
  assign _T_24066 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11}; // @[Mux.scala 19:72:@21649.4]
  assign _T_24067 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,_T_24059}; // @[Mux.scala 19:72:@21650.4]
  assign _T_24069 = _T_2692 ? _T_24067 : 16'h0; // @[Mux.scala 19:72:@21651.4]
  assign _T_24076 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@21658.4]
  assign _T_24083 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12}; // @[Mux.scala 19:72:@21665.4]
  assign _T_24084 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,_T_24076}; // @[Mux.scala 19:72:@21666.4]
  assign _T_24086 = _T_2693 ? _T_24084 : 16'h0; // @[Mux.scala 19:72:@21667.4]
  assign _T_24093 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@21674.4]
  assign _T_24100 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13}; // @[Mux.scala 19:72:@21681.4]
  assign _T_24101 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,_T_24093}; // @[Mux.scala 19:72:@21682.4]
  assign _T_24103 = _T_2694 ? _T_24101 : 16'h0; // @[Mux.scala 19:72:@21683.4]
  assign _T_24110 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@21690.4]
  assign _T_24117 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14}; // @[Mux.scala 19:72:@21697.4]
  assign _T_24118 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,_T_24110}; // @[Mux.scala 19:72:@21698.4]
  assign _T_24120 = _T_2695 ? _T_24118 : 16'h0; // @[Mux.scala 19:72:@21699.4]
  assign _T_24127 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7}; // @[Mux.scala 19:72:@21706.4]
  assign _T_24134 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15}; // @[Mux.scala 19:72:@21713.4]
  assign _T_24135 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,_T_24127}; // @[Mux.scala 19:72:@21714.4]
  assign _T_24137 = _T_2696 ? _T_24135 : 16'h0; // @[Mux.scala 19:72:@21715.4]
  assign _T_24152 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,_T_24015}; // @[Mux.scala 19:72:@21730.4]
  assign _T_24154 = _T_2697 ? _T_24152 : 16'h0; // @[Mux.scala 19:72:@21731.4]
  assign _T_24169 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,_T_24032}; // @[Mux.scala 19:72:@21746.4]
  assign _T_24171 = _T_2698 ? _T_24169 : 16'h0; // @[Mux.scala 19:72:@21747.4]
  assign _T_24186 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,_T_24049}; // @[Mux.scala 19:72:@21762.4]
  assign _T_24188 = _T_2699 ? _T_24186 : 16'h0; // @[Mux.scala 19:72:@21763.4]
  assign _T_24203 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,_T_24066}; // @[Mux.scala 19:72:@21778.4]
  assign _T_24205 = _T_2700 ? _T_24203 : 16'h0; // @[Mux.scala 19:72:@21779.4]
  assign _T_24220 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,_T_24083}; // @[Mux.scala 19:72:@21794.4]
  assign _T_24222 = _T_2701 ? _T_24220 : 16'h0; // @[Mux.scala 19:72:@21795.4]
  assign _T_24237 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,_T_24100}; // @[Mux.scala 19:72:@21810.4]
  assign _T_24239 = _T_2702 ? _T_24237 : 16'h0; // @[Mux.scala 19:72:@21811.4]
  assign _T_24254 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,_T_24117}; // @[Mux.scala 19:72:@21826.4]
  assign _T_24256 = _T_2703 ? _T_24254 : 16'h0; // @[Mux.scala 19:72:@21827.4]
  assign _T_24271 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,_T_24134}; // @[Mux.scala 19:72:@21842.4]
  assign _T_24273 = _T_2704 ? _T_24271 : 16'h0; // @[Mux.scala 19:72:@21843.4]
  assign _T_24274 = _T_24018 | _T_24035; // @[Mux.scala 19:72:@21844.4]
  assign _T_24275 = _T_24274 | _T_24052; // @[Mux.scala 19:72:@21845.4]
  assign _T_24276 = _T_24275 | _T_24069; // @[Mux.scala 19:72:@21846.4]
  assign _T_24277 = _T_24276 | _T_24086; // @[Mux.scala 19:72:@21847.4]
  assign _T_24278 = _T_24277 | _T_24103; // @[Mux.scala 19:72:@21848.4]
  assign _T_24279 = _T_24278 | _T_24120; // @[Mux.scala 19:72:@21849.4]
  assign _T_24280 = _T_24279 | _T_24137; // @[Mux.scala 19:72:@21850.4]
  assign _T_24281 = _T_24280 | _T_24154; // @[Mux.scala 19:72:@21851.4]
  assign _T_24282 = _T_24281 | _T_24171; // @[Mux.scala 19:72:@21852.4]
  assign _T_24283 = _T_24282 | _T_24188; // @[Mux.scala 19:72:@21853.4]
  assign _T_24284 = _T_24283 | _T_24205; // @[Mux.scala 19:72:@21854.4]
  assign _T_24285 = _T_24284 | _T_24222; // @[Mux.scala 19:72:@21855.4]
  assign _T_24286 = _T_24285 | _T_24239; // @[Mux.scala 19:72:@21856.4]
  assign _T_24287 = _T_24286 | _T_24256; // @[Mux.scala 19:72:@21857.4]
  assign _T_24288 = _T_24287 | _T_24273; // @[Mux.scala 19:72:@21858.4]
  assign _T_24866 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0}; // @[Mux.scala 19:72:@22208.4]
  assign _T_24873 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8}; // @[Mux.scala 19:72:@22215.4]
  assign _T_24874 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,_T_24866}; // @[Mux.scala 19:72:@22216.4]
  assign _T_24876 = _T_2689 ? _T_24874 : 16'h0; // @[Mux.scala 19:72:@22217.4]
  assign _T_24883 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1}; // @[Mux.scala 19:72:@22224.4]
  assign _T_24890 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9}; // @[Mux.scala 19:72:@22231.4]
  assign _T_24891 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,_T_24883}; // @[Mux.scala 19:72:@22232.4]
  assign _T_24893 = _T_2690 ? _T_24891 : 16'h0; // @[Mux.scala 19:72:@22233.4]
  assign _T_24900 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2}; // @[Mux.scala 19:72:@22240.4]
  assign _T_24907 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10}; // @[Mux.scala 19:72:@22247.4]
  assign _T_24908 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,_T_24900}; // @[Mux.scala 19:72:@22248.4]
  assign _T_24910 = _T_2691 ? _T_24908 : 16'h0; // @[Mux.scala 19:72:@22249.4]
  assign _T_24917 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3}; // @[Mux.scala 19:72:@22256.4]
  assign _T_24924 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11}; // @[Mux.scala 19:72:@22263.4]
  assign _T_24925 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,_T_24917}; // @[Mux.scala 19:72:@22264.4]
  assign _T_24927 = _T_2692 ? _T_24925 : 16'h0; // @[Mux.scala 19:72:@22265.4]
  assign _T_24934 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4}; // @[Mux.scala 19:72:@22272.4]
  assign _T_24941 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12}; // @[Mux.scala 19:72:@22279.4]
  assign _T_24942 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,_T_24934}; // @[Mux.scala 19:72:@22280.4]
  assign _T_24944 = _T_2693 ? _T_24942 : 16'h0; // @[Mux.scala 19:72:@22281.4]
  assign _T_24951 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5}; // @[Mux.scala 19:72:@22288.4]
  assign _T_24958 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13}; // @[Mux.scala 19:72:@22295.4]
  assign _T_24959 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,_T_24951}; // @[Mux.scala 19:72:@22296.4]
  assign _T_24961 = _T_2694 ? _T_24959 : 16'h0; // @[Mux.scala 19:72:@22297.4]
  assign _T_24968 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6}; // @[Mux.scala 19:72:@22304.4]
  assign _T_24975 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14}; // @[Mux.scala 19:72:@22311.4]
  assign _T_24976 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,_T_24968}; // @[Mux.scala 19:72:@22312.4]
  assign _T_24978 = _T_2695 ? _T_24976 : 16'h0; // @[Mux.scala 19:72:@22313.4]
  assign _T_24985 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7}; // @[Mux.scala 19:72:@22320.4]
  assign _T_24992 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15}; // @[Mux.scala 19:72:@22327.4]
  assign _T_24993 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,_T_24985}; // @[Mux.scala 19:72:@22328.4]
  assign _T_24995 = _T_2696 ? _T_24993 : 16'h0; // @[Mux.scala 19:72:@22329.4]
  assign _T_25010 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,_T_24873}; // @[Mux.scala 19:72:@22344.4]
  assign _T_25012 = _T_2697 ? _T_25010 : 16'h0; // @[Mux.scala 19:72:@22345.4]
  assign _T_25027 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,_T_24890}; // @[Mux.scala 19:72:@22360.4]
  assign _T_25029 = _T_2698 ? _T_25027 : 16'h0; // @[Mux.scala 19:72:@22361.4]
  assign _T_25044 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,_T_24907}; // @[Mux.scala 19:72:@22376.4]
  assign _T_25046 = _T_2699 ? _T_25044 : 16'h0; // @[Mux.scala 19:72:@22377.4]
  assign _T_25061 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,_T_24924}; // @[Mux.scala 19:72:@22392.4]
  assign _T_25063 = _T_2700 ? _T_25061 : 16'h0; // @[Mux.scala 19:72:@22393.4]
  assign _T_25078 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,_T_24941}; // @[Mux.scala 19:72:@22408.4]
  assign _T_25080 = _T_2701 ? _T_25078 : 16'h0; // @[Mux.scala 19:72:@22409.4]
  assign _T_25095 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,_T_24958}; // @[Mux.scala 19:72:@22424.4]
  assign _T_25097 = _T_2702 ? _T_25095 : 16'h0; // @[Mux.scala 19:72:@22425.4]
  assign _T_25112 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,_T_24975}; // @[Mux.scala 19:72:@22440.4]
  assign _T_25114 = _T_2703 ? _T_25112 : 16'h0; // @[Mux.scala 19:72:@22441.4]
  assign _T_25129 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,_T_24992}; // @[Mux.scala 19:72:@22456.4]
  assign _T_25131 = _T_2704 ? _T_25129 : 16'h0; // @[Mux.scala 19:72:@22457.4]
  assign _T_25132 = _T_24876 | _T_24893; // @[Mux.scala 19:72:@22458.4]
  assign _T_25133 = _T_25132 | _T_24910; // @[Mux.scala 19:72:@22459.4]
  assign _T_25134 = _T_25133 | _T_24927; // @[Mux.scala 19:72:@22460.4]
  assign _T_25135 = _T_25134 | _T_24944; // @[Mux.scala 19:72:@22461.4]
  assign _T_25136 = _T_25135 | _T_24961; // @[Mux.scala 19:72:@22462.4]
  assign _T_25137 = _T_25136 | _T_24978; // @[Mux.scala 19:72:@22463.4]
  assign _T_25138 = _T_25137 | _T_24995; // @[Mux.scala 19:72:@22464.4]
  assign _T_25139 = _T_25138 | _T_25012; // @[Mux.scala 19:72:@22465.4]
  assign _T_25140 = _T_25139 | _T_25029; // @[Mux.scala 19:72:@22466.4]
  assign _T_25141 = _T_25140 | _T_25046; // @[Mux.scala 19:72:@22467.4]
  assign _T_25142 = _T_25141 | _T_25063; // @[Mux.scala 19:72:@22468.4]
  assign _T_25143 = _T_25142 | _T_25080; // @[Mux.scala 19:72:@22469.4]
  assign _T_25144 = _T_25143 | _T_25097; // @[Mux.scala 19:72:@22470.4]
  assign _T_25145 = _T_25144 | _T_25114; // @[Mux.scala 19:72:@22471.4]
  assign _T_25146 = _T_25145 | _T_25131; // @[Mux.scala 19:72:@22472.4]
  assign _T_25724 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0}; // @[Mux.scala 19:72:@22822.4]
  assign _T_25731 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8}; // @[Mux.scala 19:72:@22829.4]
  assign _T_25732 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,_T_25724}; // @[Mux.scala 19:72:@22830.4]
  assign _T_25734 = _T_2689 ? _T_25732 : 16'h0; // @[Mux.scala 19:72:@22831.4]
  assign _T_25741 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1}; // @[Mux.scala 19:72:@22838.4]
  assign _T_25748 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9}; // @[Mux.scala 19:72:@22845.4]
  assign _T_25749 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,_T_25741}; // @[Mux.scala 19:72:@22846.4]
  assign _T_25751 = _T_2690 ? _T_25749 : 16'h0; // @[Mux.scala 19:72:@22847.4]
  assign _T_25758 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2}; // @[Mux.scala 19:72:@22854.4]
  assign _T_25765 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10}; // @[Mux.scala 19:72:@22861.4]
  assign _T_25766 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,_T_25758}; // @[Mux.scala 19:72:@22862.4]
  assign _T_25768 = _T_2691 ? _T_25766 : 16'h0; // @[Mux.scala 19:72:@22863.4]
  assign _T_25775 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3}; // @[Mux.scala 19:72:@22870.4]
  assign _T_25782 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11}; // @[Mux.scala 19:72:@22877.4]
  assign _T_25783 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,_T_25775}; // @[Mux.scala 19:72:@22878.4]
  assign _T_25785 = _T_2692 ? _T_25783 : 16'h0; // @[Mux.scala 19:72:@22879.4]
  assign _T_25792 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4}; // @[Mux.scala 19:72:@22886.4]
  assign _T_25799 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12}; // @[Mux.scala 19:72:@22893.4]
  assign _T_25800 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,_T_25792}; // @[Mux.scala 19:72:@22894.4]
  assign _T_25802 = _T_2693 ? _T_25800 : 16'h0; // @[Mux.scala 19:72:@22895.4]
  assign _T_25809 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5}; // @[Mux.scala 19:72:@22902.4]
  assign _T_25816 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13}; // @[Mux.scala 19:72:@22909.4]
  assign _T_25817 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,_T_25809}; // @[Mux.scala 19:72:@22910.4]
  assign _T_25819 = _T_2694 ? _T_25817 : 16'h0; // @[Mux.scala 19:72:@22911.4]
  assign _T_25826 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6}; // @[Mux.scala 19:72:@22918.4]
  assign _T_25833 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14}; // @[Mux.scala 19:72:@22925.4]
  assign _T_25834 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,_T_25826}; // @[Mux.scala 19:72:@22926.4]
  assign _T_25836 = _T_2695 ? _T_25834 : 16'h0; // @[Mux.scala 19:72:@22927.4]
  assign _T_25843 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7}; // @[Mux.scala 19:72:@22934.4]
  assign _T_25850 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15}; // @[Mux.scala 19:72:@22941.4]
  assign _T_25851 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,_T_25843}; // @[Mux.scala 19:72:@22942.4]
  assign _T_25853 = _T_2696 ? _T_25851 : 16'h0; // @[Mux.scala 19:72:@22943.4]
  assign _T_25868 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,_T_25731}; // @[Mux.scala 19:72:@22958.4]
  assign _T_25870 = _T_2697 ? _T_25868 : 16'h0; // @[Mux.scala 19:72:@22959.4]
  assign _T_25885 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,_T_25748}; // @[Mux.scala 19:72:@22974.4]
  assign _T_25887 = _T_2698 ? _T_25885 : 16'h0; // @[Mux.scala 19:72:@22975.4]
  assign _T_25902 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,_T_25765}; // @[Mux.scala 19:72:@22990.4]
  assign _T_25904 = _T_2699 ? _T_25902 : 16'h0; // @[Mux.scala 19:72:@22991.4]
  assign _T_25919 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,_T_25782}; // @[Mux.scala 19:72:@23006.4]
  assign _T_25921 = _T_2700 ? _T_25919 : 16'h0; // @[Mux.scala 19:72:@23007.4]
  assign _T_25936 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,_T_25799}; // @[Mux.scala 19:72:@23022.4]
  assign _T_25938 = _T_2701 ? _T_25936 : 16'h0; // @[Mux.scala 19:72:@23023.4]
  assign _T_25953 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,_T_25816}; // @[Mux.scala 19:72:@23038.4]
  assign _T_25955 = _T_2702 ? _T_25953 : 16'h0; // @[Mux.scala 19:72:@23039.4]
  assign _T_25970 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,_T_25833}; // @[Mux.scala 19:72:@23054.4]
  assign _T_25972 = _T_2703 ? _T_25970 : 16'h0; // @[Mux.scala 19:72:@23055.4]
  assign _T_25987 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,_T_25850}; // @[Mux.scala 19:72:@23070.4]
  assign _T_25989 = _T_2704 ? _T_25987 : 16'h0; // @[Mux.scala 19:72:@23071.4]
  assign _T_25990 = _T_25734 | _T_25751; // @[Mux.scala 19:72:@23072.4]
  assign _T_25991 = _T_25990 | _T_25768; // @[Mux.scala 19:72:@23073.4]
  assign _T_25992 = _T_25991 | _T_25785; // @[Mux.scala 19:72:@23074.4]
  assign _T_25993 = _T_25992 | _T_25802; // @[Mux.scala 19:72:@23075.4]
  assign _T_25994 = _T_25993 | _T_25819; // @[Mux.scala 19:72:@23076.4]
  assign _T_25995 = _T_25994 | _T_25836; // @[Mux.scala 19:72:@23077.4]
  assign _T_25996 = _T_25995 | _T_25853; // @[Mux.scala 19:72:@23078.4]
  assign _T_25997 = _T_25996 | _T_25870; // @[Mux.scala 19:72:@23079.4]
  assign _T_25998 = _T_25997 | _T_25887; // @[Mux.scala 19:72:@23080.4]
  assign _T_25999 = _T_25998 | _T_25904; // @[Mux.scala 19:72:@23081.4]
  assign _T_26000 = _T_25999 | _T_25921; // @[Mux.scala 19:72:@23082.4]
  assign _T_26001 = _T_26000 | _T_25938; // @[Mux.scala 19:72:@23083.4]
  assign _T_26002 = _T_26001 | _T_25955; // @[Mux.scala 19:72:@23084.4]
  assign _T_26003 = _T_26002 | _T_25972; // @[Mux.scala 19:72:@23085.4]
  assign _T_26004 = _T_26003 | _T_25989; // @[Mux.scala 19:72:@23086.4]
  assign _T_26582 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0}; // @[Mux.scala 19:72:@23436.4]
  assign _T_26589 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8}; // @[Mux.scala 19:72:@23443.4]
  assign _T_26590 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,_T_26582}; // @[Mux.scala 19:72:@23444.4]
  assign _T_26592 = _T_2689 ? _T_26590 : 16'h0; // @[Mux.scala 19:72:@23445.4]
  assign _T_26599 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1}; // @[Mux.scala 19:72:@23452.4]
  assign _T_26606 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9}; // @[Mux.scala 19:72:@23459.4]
  assign _T_26607 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,_T_26599}; // @[Mux.scala 19:72:@23460.4]
  assign _T_26609 = _T_2690 ? _T_26607 : 16'h0; // @[Mux.scala 19:72:@23461.4]
  assign _T_26616 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2}; // @[Mux.scala 19:72:@23468.4]
  assign _T_26623 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10}; // @[Mux.scala 19:72:@23475.4]
  assign _T_26624 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,_T_26616}; // @[Mux.scala 19:72:@23476.4]
  assign _T_26626 = _T_2691 ? _T_26624 : 16'h0; // @[Mux.scala 19:72:@23477.4]
  assign _T_26633 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3}; // @[Mux.scala 19:72:@23484.4]
  assign _T_26640 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11}; // @[Mux.scala 19:72:@23491.4]
  assign _T_26641 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,_T_26633}; // @[Mux.scala 19:72:@23492.4]
  assign _T_26643 = _T_2692 ? _T_26641 : 16'h0; // @[Mux.scala 19:72:@23493.4]
  assign _T_26650 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4}; // @[Mux.scala 19:72:@23500.4]
  assign _T_26657 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12}; // @[Mux.scala 19:72:@23507.4]
  assign _T_26658 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,_T_26650}; // @[Mux.scala 19:72:@23508.4]
  assign _T_26660 = _T_2693 ? _T_26658 : 16'h0; // @[Mux.scala 19:72:@23509.4]
  assign _T_26667 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5}; // @[Mux.scala 19:72:@23516.4]
  assign _T_26674 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13}; // @[Mux.scala 19:72:@23523.4]
  assign _T_26675 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,_T_26667}; // @[Mux.scala 19:72:@23524.4]
  assign _T_26677 = _T_2694 ? _T_26675 : 16'h0; // @[Mux.scala 19:72:@23525.4]
  assign _T_26684 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6}; // @[Mux.scala 19:72:@23532.4]
  assign _T_26691 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14}; // @[Mux.scala 19:72:@23539.4]
  assign _T_26692 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,_T_26684}; // @[Mux.scala 19:72:@23540.4]
  assign _T_26694 = _T_2695 ? _T_26692 : 16'h0; // @[Mux.scala 19:72:@23541.4]
  assign _T_26701 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7}; // @[Mux.scala 19:72:@23548.4]
  assign _T_26708 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15}; // @[Mux.scala 19:72:@23555.4]
  assign _T_26709 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,_T_26701}; // @[Mux.scala 19:72:@23556.4]
  assign _T_26711 = _T_2696 ? _T_26709 : 16'h0; // @[Mux.scala 19:72:@23557.4]
  assign _T_26726 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,_T_26589}; // @[Mux.scala 19:72:@23572.4]
  assign _T_26728 = _T_2697 ? _T_26726 : 16'h0; // @[Mux.scala 19:72:@23573.4]
  assign _T_26743 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,_T_26606}; // @[Mux.scala 19:72:@23588.4]
  assign _T_26745 = _T_2698 ? _T_26743 : 16'h0; // @[Mux.scala 19:72:@23589.4]
  assign _T_26760 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,_T_26623}; // @[Mux.scala 19:72:@23604.4]
  assign _T_26762 = _T_2699 ? _T_26760 : 16'h0; // @[Mux.scala 19:72:@23605.4]
  assign _T_26777 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,_T_26640}; // @[Mux.scala 19:72:@23620.4]
  assign _T_26779 = _T_2700 ? _T_26777 : 16'h0; // @[Mux.scala 19:72:@23621.4]
  assign _T_26794 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,_T_26657}; // @[Mux.scala 19:72:@23636.4]
  assign _T_26796 = _T_2701 ? _T_26794 : 16'h0; // @[Mux.scala 19:72:@23637.4]
  assign _T_26811 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,_T_26674}; // @[Mux.scala 19:72:@23652.4]
  assign _T_26813 = _T_2702 ? _T_26811 : 16'h0; // @[Mux.scala 19:72:@23653.4]
  assign _T_26828 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,_T_26691}; // @[Mux.scala 19:72:@23668.4]
  assign _T_26830 = _T_2703 ? _T_26828 : 16'h0; // @[Mux.scala 19:72:@23669.4]
  assign _T_26845 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,_T_26708}; // @[Mux.scala 19:72:@23684.4]
  assign _T_26847 = _T_2704 ? _T_26845 : 16'h0; // @[Mux.scala 19:72:@23685.4]
  assign _T_26848 = _T_26592 | _T_26609; // @[Mux.scala 19:72:@23686.4]
  assign _T_26849 = _T_26848 | _T_26626; // @[Mux.scala 19:72:@23687.4]
  assign _T_26850 = _T_26849 | _T_26643; // @[Mux.scala 19:72:@23688.4]
  assign _T_26851 = _T_26850 | _T_26660; // @[Mux.scala 19:72:@23689.4]
  assign _T_26852 = _T_26851 | _T_26677; // @[Mux.scala 19:72:@23690.4]
  assign _T_26853 = _T_26852 | _T_26694; // @[Mux.scala 19:72:@23691.4]
  assign _T_26854 = _T_26853 | _T_26711; // @[Mux.scala 19:72:@23692.4]
  assign _T_26855 = _T_26854 | _T_26728; // @[Mux.scala 19:72:@23693.4]
  assign _T_26856 = _T_26855 | _T_26745; // @[Mux.scala 19:72:@23694.4]
  assign _T_26857 = _T_26856 | _T_26762; // @[Mux.scala 19:72:@23695.4]
  assign _T_26858 = _T_26857 | _T_26779; // @[Mux.scala 19:72:@23696.4]
  assign _T_26859 = _T_26858 | _T_26796; // @[Mux.scala 19:72:@23697.4]
  assign _T_26860 = _T_26859 | _T_26813; // @[Mux.scala 19:72:@23698.4]
  assign _T_26861 = _T_26860 | _T_26830; // @[Mux.scala 19:72:@23699.4]
  assign _T_26862 = _T_26861 | _T_26847; // @[Mux.scala 19:72:@23700.4]
  assign _T_27440 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0}; // @[Mux.scala 19:72:@24050.4]
  assign _T_27447 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8}; // @[Mux.scala 19:72:@24057.4]
  assign _T_27448 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,_T_27440}; // @[Mux.scala 19:72:@24058.4]
  assign _T_27450 = _T_2689 ? _T_27448 : 16'h0; // @[Mux.scala 19:72:@24059.4]
  assign _T_27457 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1}; // @[Mux.scala 19:72:@24066.4]
  assign _T_27464 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9}; // @[Mux.scala 19:72:@24073.4]
  assign _T_27465 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,_T_27457}; // @[Mux.scala 19:72:@24074.4]
  assign _T_27467 = _T_2690 ? _T_27465 : 16'h0; // @[Mux.scala 19:72:@24075.4]
  assign _T_27474 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2}; // @[Mux.scala 19:72:@24082.4]
  assign _T_27481 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10}; // @[Mux.scala 19:72:@24089.4]
  assign _T_27482 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,_T_27474}; // @[Mux.scala 19:72:@24090.4]
  assign _T_27484 = _T_2691 ? _T_27482 : 16'h0; // @[Mux.scala 19:72:@24091.4]
  assign _T_27491 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3}; // @[Mux.scala 19:72:@24098.4]
  assign _T_27498 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11}; // @[Mux.scala 19:72:@24105.4]
  assign _T_27499 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,_T_27491}; // @[Mux.scala 19:72:@24106.4]
  assign _T_27501 = _T_2692 ? _T_27499 : 16'h0; // @[Mux.scala 19:72:@24107.4]
  assign _T_27508 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4}; // @[Mux.scala 19:72:@24114.4]
  assign _T_27515 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12}; // @[Mux.scala 19:72:@24121.4]
  assign _T_27516 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,_T_27508}; // @[Mux.scala 19:72:@24122.4]
  assign _T_27518 = _T_2693 ? _T_27516 : 16'h0; // @[Mux.scala 19:72:@24123.4]
  assign _T_27525 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5}; // @[Mux.scala 19:72:@24130.4]
  assign _T_27532 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13}; // @[Mux.scala 19:72:@24137.4]
  assign _T_27533 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,_T_27525}; // @[Mux.scala 19:72:@24138.4]
  assign _T_27535 = _T_2694 ? _T_27533 : 16'h0; // @[Mux.scala 19:72:@24139.4]
  assign _T_27542 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6}; // @[Mux.scala 19:72:@24146.4]
  assign _T_27549 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14}; // @[Mux.scala 19:72:@24153.4]
  assign _T_27550 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,_T_27542}; // @[Mux.scala 19:72:@24154.4]
  assign _T_27552 = _T_2695 ? _T_27550 : 16'h0; // @[Mux.scala 19:72:@24155.4]
  assign _T_27559 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7}; // @[Mux.scala 19:72:@24162.4]
  assign _T_27566 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15}; // @[Mux.scala 19:72:@24169.4]
  assign _T_27567 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,_T_27559}; // @[Mux.scala 19:72:@24170.4]
  assign _T_27569 = _T_2696 ? _T_27567 : 16'h0; // @[Mux.scala 19:72:@24171.4]
  assign _T_27584 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,_T_27447}; // @[Mux.scala 19:72:@24186.4]
  assign _T_27586 = _T_2697 ? _T_27584 : 16'h0; // @[Mux.scala 19:72:@24187.4]
  assign _T_27601 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,_T_27464}; // @[Mux.scala 19:72:@24202.4]
  assign _T_27603 = _T_2698 ? _T_27601 : 16'h0; // @[Mux.scala 19:72:@24203.4]
  assign _T_27618 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,_T_27481}; // @[Mux.scala 19:72:@24218.4]
  assign _T_27620 = _T_2699 ? _T_27618 : 16'h0; // @[Mux.scala 19:72:@24219.4]
  assign _T_27635 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,_T_27498}; // @[Mux.scala 19:72:@24234.4]
  assign _T_27637 = _T_2700 ? _T_27635 : 16'h0; // @[Mux.scala 19:72:@24235.4]
  assign _T_27652 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,_T_27515}; // @[Mux.scala 19:72:@24250.4]
  assign _T_27654 = _T_2701 ? _T_27652 : 16'h0; // @[Mux.scala 19:72:@24251.4]
  assign _T_27669 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,_T_27532}; // @[Mux.scala 19:72:@24266.4]
  assign _T_27671 = _T_2702 ? _T_27669 : 16'h0; // @[Mux.scala 19:72:@24267.4]
  assign _T_27686 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,_T_27549}; // @[Mux.scala 19:72:@24282.4]
  assign _T_27688 = _T_2703 ? _T_27686 : 16'h0; // @[Mux.scala 19:72:@24283.4]
  assign _T_27703 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,_T_27566}; // @[Mux.scala 19:72:@24298.4]
  assign _T_27705 = _T_2704 ? _T_27703 : 16'h0; // @[Mux.scala 19:72:@24299.4]
  assign _T_27706 = _T_27450 | _T_27467; // @[Mux.scala 19:72:@24300.4]
  assign _T_27707 = _T_27706 | _T_27484; // @[Mux.scala 19:72:@24301.4]
  assign _T_27708 = _T_27707 | _T_27501; // @[Mux.scala 19:72:@24302.4]
  assign _T_27709 = _T_27708 | _T_27518; // @[Mux.scala 19:72:@24303.4]
  assign _T_27710 = _T_27709 | _T_27535; // @[Mux.scala 19:72:@24304.4]
  assign _T_27711 = _T_27710 | _T_27552; // @[Mux.scala 19:72:@24305.4]
  assign _T_27712 = _T_27711 | _T_27569; // @[Mux.scala 19:72:@24306.4]
  assign _T_27713 = _T_27712 | _T_27586; // @[Mux.scala 19:72:@24307.4]
  assign _T_27714 = _T_27713 | _T_27603; // @[Mux.scala 19:72:@24308.4]
  assign _T_27715 = _T_27714 | _T_27620; // @[Mux.scala 19:72:@24309.4]
  assign _T_27716 = _T_27715 | _T_27637; // @[Mux.scala 19:72:@24310.4]
  assign _T_27717 = _T_27716 | _T_27654; // @[Mux.scala 19:72:@24311.4]
  assign _T_27718 = _T_27717 | _T_27671; // @[Mux.scala 19:72:@24312.4]
  assign _T_27719 = _T_27718 | _T_27688; // @[Mux.scala 19:72:@24313.4]
  assign _T_27720 = _T_27719 | _T_27705; // @[Mux.scala 19:72:@24314.4]
  assign _T_28298 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0}; // @[Mux.scala 19:72:@24664.4]
  assign _T_28305 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8}; // @[Mux.scala 19:72:@24671.4]
  assign _T_28306 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,_T_28298}; // @[Mux.scala 19:72:@24672.4]
  assign _T_28308 = _T_2689 ? _T_28306 : 16'h0; // @[Mux.scala 19:72:@24673.4]
  assign _T_28315 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1}; // @[Mux.scala 19:72:@24680.4]
  assign _T_28322 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9}; // @[Mux.scala 19:72:@24687.4]
  assign _T_28323 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,_T_28315}; // @[Mux.scala 19:72:@24688.4]
  assign _T_28325 = _T_2690 ? _T_28323 : 16'h0; // @[Mux.scala 19:72:@24689.4]
  assign _T_28332 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2}; // @[Mux.scala 19:72:@24696.4]
  assign _T_28339 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10}; // @[Mux.scala 19:72:@24703.4]
  assign _T_28340 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,_T_28332}; // @[Mux.scala 19:72:@24704.4]
  assign _T_28342 = _T_2691 ? _T_28340 : 16'h0; // @[Mux.scala 19:72:@24705.4]
  assign _T_28349 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3}; // @[Mux.scala 19:72:@24712.4]
  assign _T_28356 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11}; // @[Mux.scala 19:72:@24719.4]
  assign _T_28357 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,_T_28349}; // @[Mux.scala 19:72:@24720.4]
  assign _T_28359 = _T_2692 ? _T_28357 : 16'h0; // @[Mux.scala 19:72:@24721.4]
  assign _T_28366 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4}; // @[Mux.scala 19:72:@24728.4]
  assign _T_28373 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12}; // @[Mux.scala 19:72:@24735.4]
  assign _T_28374 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,_T_28366}; // @[Mux.scala 19:72:@24736.4]
  assign _T_28376 = _T_2693 ? _T_28374 : 16'h0; // @[Mux.scala 19:72:@24737.4]
  assign _T_28383 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5}; // @[Mux.scala 19:72:@24744.4]
  assign _T_28390 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13}; // @[Mux.scala 19:72:@24751.4]
  assign _T_28391 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,_T_28383}; // @[Mux.scala 19:72:@24752.4]
  assign _T_28393 = _T_2694 ? _T_28391 : 16'h0; // @[Mux.scala 19:72:@24753.4]
  assign _T_28400 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6}; // @[Mux.scala 19:72:@24760.4]
  assign _T_28407 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14}; // @[Mux.scala 19:72:@24767.4]
  assign _T_28408 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,_T_28400}; // @[Mux.scala 19:72:@24768.4]
  assign _T_28410 = _T_2695 ? _T_28408 : 16'h0; // @[Mux.scala 19:72:@24769.4]
  assign _T_28417 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7}; // @[Mux.scala 19:72:@24776.4]
  assign _T_28424 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15}; // @[Mux.scala 19:72:@24783.4]
  assign _T_28425 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,_T_28417}; // @[Mux.scala 19:72:@24784.4]
  assign _T_28427 = _T_2696 ? _T_28425 : 16'h0; // @[Mux.scala 19:72:@24785.4]
  assign _T_28442 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,_T_28305}; // @[Mux.scala 19:72:@24800.4]
  assign _T_28444 = _T_2697 ? _T_28442 : 16'h0; // @[Mux.scala 19:72:@24801.4]
  assign _T_28459 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,_T_28322}; // @[Mux.scala 19:72:@24816.4]
  assign _T_28461 = _T_2698 ? _T_28459 : 16'h0; // @[Mux.scala 19:72:@24817.4]
  assign _T_28476 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,_T_28339}; // @[Mux.scala 19:72:@24832.4]
  assign _T_28478 = _T_2699 ? _T_28476 : 16'h0; // @[Mux.scala 19:72:@24833.4]
  assign _T_28493 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,_T_28356}; // @[Mux.scala 19:72:@24848.4]
  assign _T_28495 = _T_2700 ? _T_28493 : 16'h0; // @[Mux.scala 19:72:@24849.4]
  assign _T_28510 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,_T_28373}; // @[Mux.scala 19:72:@24864.4]
  assign _T_28512 = _T_2701 ? _T_28510 : 16'h0; // @[Mux.scala 19:72:@24865.4]
  assign _T_28527 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,_T_28390}; // @[Mux.scala 19:72:@24880.4]
  assign _T_28529 = _T_2702 ? _T_28527 : 16'h0; // @[Mux.scala 19:72:@24881.4]
  assign _T_28544 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,_T_28407}; // @[Mux.scala 19:72:@24896.4]
  assign _T_28546 = _T_2703 ? _T_28544 : 16'h0; // @[Mux.scala 19:72:@24897.4]
  assign _T_28561 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,_T_28424}; // @[Mux.scala 19:72:@24912.4]
  assign _T_28563 = _T_2704 ? _T_28561 : 16'h0; // @[Mux.scala 19:72:@24913.4]
  assign _T_28564 = _T_28308 | _T_28325; // @[Mux.scala 19:72:@24914.4]
  assign _T_28565 = _T_28564 | _T_28342; // @[Mux.scala 19:72:@24915.4]
  assign _T_28566 = _T_28565 | _T_28359; // @[Mux.scala 19:72:@24916.4]
  assign _T_28567 = _T_28566 | _T_28376; // @[Mux.scala 19:72:@24917.4]
  assign _T_28568 = _T_28567 | _T_28393; // @[Mux.scala 19:72:@24918.4]
  assign _T_28569 = _T_28568 | _T_28410; // @[Mux.scala 19:72:@24919.4]
  assign _T_28570 = _T_28569 | _T_28427; // @[Mux.scala 19:72:@24920.4]
  assign _T_28571 = _T_28570 | _T_28444; // @[Mux.scala 19:72:@24921.4]
  assign _T_28572 = _T_28571 | _T_28461; // @[Mux.scala 19:72:@24922.4]
  assign _T_28573 = _T_28572 | _T_28478; // @[Mux.scala 19:72:@24923.4]
  assign _T_28574 = _T_28573 | _T_28495; // @[Mux.scala 19:72:@24924.4]
  assign _T_28575 = _T_28574 | _T_28512; // @[Mux.scala 19:72:@24925.4]
  assign _T_28576 = _T_28575 | _T_28529; // @[Mux.scala 19:72:@24926.4]
  assign _T_28577 = _T_28576 | _T_28546; // @[Mux.scala 19:72:@24927.4]
  assign _T_28578 = _T_28577 | _T_28563; // @[Mux.scala 19:72:@24928.4]
  assign _T_29156 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0}; // @[Mux.scala 19:72:@25278.4]
  assign _T_29163 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8}; // @[Mux.scala 19:72:@25285.4]
  assign _T_29164 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,_T_29156}; // @[Mux.scala 19:72:@25286.4]
  assign _T_29166 = _T_2689 ? _T_29164 : 16'h0; // @[Mux.scala 19:72:@25287.4]
  assign _T_29173 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1}; // @[Mux.scala 19:72:@25294.4]
  assign _T_29180 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9}; // @[Mux.scala 19:72:@25301.4]
  assign _T_29181 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,_T_29173}; // @[Mux.scala 19:72:@25302.4]
  assign _T_29183 = _T_2690 ? _T_29181 : 16'h0; // @[Mux.scala 19:72:@25303.4]
  assign _T_29190 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2}; // @[Mux.scala 19:72:@25310.4]
  assign _T_29197 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10}; // @[Mux.scala 19:72:@25317.4]
  assign _T_29198 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,_T_29190}; // @[Mux.scala 19:72:@25318.4]
  assign _T_29200 = _T_2691 ? _T_29198 : 16'h0; // @[Mux.scala 19:72:@25319.4]
  assign _T_29207 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3}; // @[Mux.scala 19:72:@25326.4]
  assign _T_29214 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11}; // @[Mux.scala 19:72:@25333.4]
  assign _T_29215 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,_T_29207}; // @[Mux.scala 19:72:@25334.4]
  assign _T_29217 = _T_2692 ? _T_29215 : 16'h0; // @[Mux.scala 19:72:@25335.4]
  assign _T_29224 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4}; // @[Mux.scala 19:72:@25342.4]
  assign _T_29231 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12}; // @[Mux.scala 19:72:@25349.4]
  assign _T_29232 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,_T_29224}; // @[Mux.scala 19:72:@25350.4]
  assign _T_29234 = _T_2693 ? _T_29232 : 16'h0; // @[Mux.scala 19:72:@25351.4]
  assign _T_29241 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5}; // @[Mux.scala 19:72:@25358.4]
  assign _T_29248 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13}; // @[Mux.scala 19:72:@25365.4]
  assign _T_29249 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,_T_29241}; // @[Mux.scala 19:72:@25366.4]
  assign _T_29251 = _T_2694 ? _T_29249 : 16'h0; // @[Mux.scala 19:72:@25367.4]
  assign _T_29258 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6}; // @[Mux.scala 19:72:@25374.4]
  assign _T_29265 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14}; // @[Mux.scala 19:72:@25381.4]
  assign _T_29266 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,_T_29258}; // @[Mux.scala 19:72:@25382.4]
  assign _T_29268 = _T_2695 ? _T_29266 : 16'h0; // @[Mux.scala 19:72:@25383.4]
  assign _T_29275 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7}; // @[Mux.scala 19:72:@25390.4]
  assign _T_29282 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15}; // @[Mux.scala 19:72:@25397.4]
  assign _T_29283 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,_T_29275}; // @[Mux.scala 19:72:@25398.4]
  assign _T_29285 = _T_2696 ? _T_29283 : 16'h0; // @[Mux.scala 19:72:@25399.4]
  assign _T_29300 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,_T_29163}; // @[Mux.scala 19:72:@25414.4]
  assign _T_29302 = _T_2697 ? _T_29300 : 16'h0; // @[Mux.scala 19:72:@25415.4]
  assign _T_29317 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,_T_29180}; // @[Mux.scala 19:72:@25430.4]
  assign _T_29319 = _T_2698 ? _T_29317 : 16'h0; // @[Mux.scala 19:72:@25431.4]
  assign _T_29334 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,_T_29197}; // @[Mux.scala 19:72:@25446.4]
  assign _T_29336 = _T_2699 ? _T_29334 : 16'h0; // @[Mux.scala 19:72:@25447.4]
  assign _T_29351 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,_T_29214}; // @[Mux.scala 19:72:@25462.4]
  assign _T_29353 = _T_2700 ? _T_29351 : 16'h0; // @[Mux.scala 19:72:@25463.4]
  assign _T_29368 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,_T_29231}; // @[Mux.scala 19:72:@25478.4]
  assign _T_29370 = _T_2701 ? _T_29368 : 16'h0; // @[Mux.scala 19:72:@25479.4]
  assign _T_29385 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,_T_29248}; // @[Mux.scala 19:72:@25494.4]
  assign _T_29387 = _T_2702 ? _T_29385 : 16'h0; // @[Mux.scala 19:72:@25495.4]
  assign _T_29402 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,_T_29265}; // @[Mux.scala 19:72:@25510.4]
  assign _T_29404 = _T_2703 ? _T_29402 : 16'h0; // @[Mux.scala 19:72:@25511.4]
  assign _T_29419 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,_T_29282}; // @[Mux.scala 19:72:@25526.4]
  assign _T_29421 = _T_2704 ? _T_29419 : 16'h0; // @[Mux.scala 19:72:@25527.4]
  assign _T_29422 = _T_29166 | _T_29183; // @[Mux.scala 19:72:@25528.4]
  assign _T_29423 = _T_29422 | _T_29200; // @[Mux.scala 19:72:@25529.4]
  assign _T_29424 = _T_29423 | _T_29217; // @[Mux.scala 19:72:@25530.4]
  assign _T_29425 = _T_29424 | _T_29234; // @[Mux.scala 19:72:@25531.4]
  assign _T_29426 = _T_29425 | _T_29251; // @[Mux.scala 19:72:@25532.4]
  assign _T_29427 = _T_29426 | _T_29268; // @[Mux.scala 19:72:@25533.4]
  assign _T_29428 = _T_29427 | _T_29285; // @[Mux.scala 19:72:@25534.4]
  assign _T_29429 = _T_29428 | _T_29302; // @[Mux.scala 19:72:@25535.4]
  assign _T_29430 = _T_29429 | _T_29319; // @[Mux.scala 19:72:@25536.4]
  assign _T_29431 = _T_29430 | _T_29336; // @[Mux.scala 19:72:@25537.4]
  assign _T_29432 = _T_29431 | _T_29353; // @[Mux.scala 19:72:@25538.4]
  assign _T_29433 = _T_29432 | _T_29370; // @[Mux.scala 19:72:@25539.4]
  assign _T_29434 = _T_29433 | _T_29387; // @[Mux.scala 19:72:@25540.4]
  assign _T_29435 = _T_29434 | _T_29404; // @[Mux.scala 19:72:@25541.4]
  assign _T_29436 = _T_29435 | _T_29421; // @[Mux.scala 19:72:@25542.4]
  assign _T_30014 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0}; // @[Mux.scala 19:72:@25892.4]
  assign _T_30021 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8}; // @[Mux.scala 19:72:@25899.4]
  assign _T_30022 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,_T_30014}; // @[Mux.scala 19:72:@25900.4]
  assign _T_30024 = _T_2689 ? _T_30022 : 16'h0; // @[Mux.scala 19:72:@25901.4]
  assign _T_30031 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1}; // @[Mux.scala 19:72:@25908.4]
  assign _T_30038 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9}; // @[Mux.scala 19:72:@25915.4]
  assign _T_30039 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,_T_30031}; // @[Mux.scala 19:72:@25916.4]
  assign _T_30041 = _T_2690 ? _T_30039 : 16'h0; // @[Mux.scala 19:72:@25917.4]
  assign _T_30048 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2}; // @[Mux.scala 19:72:@25924.4]
  assign _T_30055 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10}; // @[Mux.scala 19:72:@25931.4]
  assign _T_30056 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,_T_30048}; // @[Mux.scala 19:72:@25932.4]
  assign _T_30058 = _T_2691 ? _T_30056 : 16'h0; // @[Mux.scala 19:72:@25933.4]
  assign _T_30065 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3}; // @[Mux.scala 19:72:@25940.4]
  assign _T_30072 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11}; // @[Mux.scala 19:72:@25947.4]
  assign _T_30073 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,_T_30065}; // @[Mux.scala 19:72:@25948.4]
  assign _T_30075 = _T_2692 ? _T_30073 : 16'h0; // @[Mux.scala 19:72:@25949.4]
  assign _T_30082 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4}; // @[Mux.scala 19:72:@25956.4]
  assign _T_30089 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12}; // @[Mux.scala 19:72:@25963.4]
  assign _T_30090 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,_T_30082}; // @[Mux.scala 19:72:@25964.4]
  assign _T_30092 = _T_2693 ? _T_30090 : 16'h0; // @[Mux.scala 19:72:@25965.4]
  assign _T_30099 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5}; // @[Mux.scala 19:72:@25972.4]
  assign _T_30106 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13}; // @[Mux.scala 19:72:@25979.4]
  assign _T_30107 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,_T_30099}; // @[Mux.scala 19:72:@25980.4]
  assign _T_30109 = _T_2694 ? _T_30107 : 16'h0; // @[Mux.scala 19:72:@25981.4]
  assign _T_30116 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6}; // @[Mux.scala 19:72:@25988.4]
  assign _T_30123 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14}; // @[Mux.scala 19:72:@25995.4]
  assign _T_30124 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,_T_30116}; // @[Mux.scala 19:72:@25996.4]
  assign _T_30126 = _T_2695 ? _T_30124 : 16'h0; // @[Mux.scala 19:72:@25997.4]
  assign _T_30133 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7}; // @[Mux.scala 19:72:@26004.4]
  assign _T_30140 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15}; // @[Mux.scala 19:72:@26011.4]
  assign _T_30141 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,_T_30133}; // @[Mux.scala 19:72:@26012.4]
  assign _T_30143 = _T_2696 ? _T_30141 : 16'h0; // @[Mux.scala 19:72:@26013.4]
  assign _T_30158 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,_T_30021}; // @[Mux.scala 19:72:@26028.4]
  assign _T_30160 = _T_2697 ? _T_30158 : 16'h0; // @[Mux.scala 19:72:@26029.4]
  assign _T_30175 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,_T_30038}; // @[Mux.scala 19:72:@26044.4]
  assign _T_30177 = _T_2698 ? _T_30175 : 16'h0; // @[Mux.scala 19:72:@26045.4]
  assign _T_30192 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,_T_30055}; // @[Mux.scala 19:72:@26060.4]
  assign _T_30194 = _T_2699 ? _T_30192 : 16'h0; // @[Mux.scala 19:72:@26061.4]
  assign _T_30209 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,_T_30072}; // @[Mux.scala 19:72:@26076.4]
  assign _T_30211 = _T_2700 ? _T_30209 : 16'h0; // @[Mux.scala 19:72:@26077.4]
  assign _T_30226 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,_T_30089}; // @[Mux.scala 19:72:@26092.4]
  assign _T_30228 = _T_2701 ? _T_30226 : 16'h0; // @[Mux.scala 19:72:@26093.4]
  assign _T_30243 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,_T_30106}; // @[Mux.scala 19:72:@26108.4]
  assign _T_30245 = _T_2702 ? _T_30243 : 16'h0; // @[Mux.scala 19:72:@26109.4]
  assign _T_30260 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,_T_30123}; // @[Mux.scala 19:72:@26124.4]
  assign _T_30262 = _T_2703 ? _T_30260 : 16'h0; // @[Mux.scala 19:72:@26125.4]
  assign _T_30277 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,_T_30140}; // @[Mux.scala 19:72:@26140.4]
  assign _T_30279 = _T_2704 ? _T_30277 : 16'h0; // @[Mux.scala 19:72:@26141.4]
  assign _T_30280 = _T_30024 | _T_30041; // @[Mux.scala 19:72:@26142.4]
  assign _T_30281 = _T_30280 | _T_30058; // @[Mux.scala 19:72:@26143.4]
  assign _T_30282 = _T_30281 | _T_30075; // @[Mux.scala 19:72:@26144.4]
  assign _T_30283 = _T_30282 | _T_30092; // @[Mux.scala 19:72:@26145.4]
  assign _T_30284 = _T_30283 | _T_30109; // @[Mux.scala 19:72:@26146.4]
  assign _T_30285 = _T_30284 | _T_30126; // @[Mux.scala 19:72:@26147.4]
  assign _T_30286 = _T_30285 | _T_30143; // @[Mux.scala 19:72:@26148.4]
  assign _T_30287 = _T_30286 | _T_30160; // @[Mux.scala 19:72:@26149.4]
  assign _T_30288 = _T_30287 | _T_30177; // @[Mux.scala 19:72:@26150.4]
  assign _T_30289 = _T_30288 | _T_30194; // @[Mux.scala 19:72:@26151.4]
  assign _T_30290 = _T_30289 | _T_30211; // @[Mux.scala 19:72:@26152.4]
  assign _T_30291 = _T_30290 | _T_30228; // @[Mux.scala 19:72:@26153.4]
  assign _T_30292 = _T_30291 | _T_30245; // @[Mux.scala 19:72:@26154.4]
  assign _T_30293 = _T_30292 | _T_30262; // @[Mux.scala 19:72:@26155.4]
  assign _T_30294 = _T_30293 | _T_30279; // @[Mux.scala 19:72:@26156.4]
  assign _T_30872 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0}; // @[Mux.scala 19:72:@26506.4]
  assign _T_30879 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8}; // @[Mux.scala 19:72:@26513.4]
  assign _T_30880 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,_T_30872}; // @[Mux.scala 19:72:@26514.4]
  assign _T_30882 = _T_2689 ? _T_30880 : 16'h0; // @[Mux.scala 19:72:@26515.4]
  assign _T_30889 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1}; // @[Mux.scala 19:72:@26522.4]
  assign _T_30896 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9}; // @[Mux.scala 19:72:@26529.4]
  assign _T_30897 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,_T_30889}; // @[Mux.scala 19:72:@26530.4]
  assign _T_30899 = _T_2690 ? _T_30897 : 16'h0; // @[Mux.scala 19:72:@26531.4]
  assign _T_30906 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2}; // @[Mux.scala 19:72:@26538.4]
  assign _T_30913 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10}; // @[Mux.scala 19:72:@26545.4]
  assign _T_30914 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,_T_30906}; // @[Mux.scala 19:72:@26546.4]
  assign _T_30916 = _T_2691 ? _T_30914 : 16'h0; // @[Mux.scala 19:72:@26547.4]
  assign _T_30923 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3}; // @[Mux.scala 19:72:@26554.4]
  assign _T_30930 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11}; // @[Mux.scala 19:72:@26561.4]
  assign _T_30931 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,_T_30923}; // @[Mux.scala 19:72:@26562.4]
  assign _T_30933 = _T_2692 ? _T_30931 : 16'h0; // @[Mux.scala 19:72:@26563.4]
  assign _T_30940 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4}; // @[Mux.scala 19:72:@26570.4]
  assign _T_30947 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12}; // @[Mux.scala 19:72:@26577.4]
  assign _T_30948 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,_T_30940}; // @[Mux.scala 19:72:@26578.4]
  assign _T_30950 = _T_2693 ? _T_30948 : 16'h0; // @[Mux.scala 19:72:@26579.4]
  assign _T_30957 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5}; // @[Mux.scala 19:72:@26586.4]
  assign _T_30964 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13}; // @[Mux.scala 19:72:@26593.4]
  assign _T_30965 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,_T_30957}; // @[Mux.scala 19:72:@26594.4]
  assign _T_30967 = _T_2694 ? _T_30965 : 16'h0; // @[Mux.scala 19:72:@26595.4]
  assign _T_30974 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6}; // @[Mux.scala 19:72:@26602.4]
  assign _T_30981 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14}; // @[Mux.scala 19:72:@26609.4]
  assign _T_30982 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,_T_30974}; // @[Mux.scala 19:72:@26610.4]
  assign _T_30984 = _T_2695 ? _T_30982 : 16'h0; // @[Mux.scala 19:72:@26611.4]
  assign _T_30991 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7}; // @[Mux.scala 19:72:@26618.4]
  assign _T_30998 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15}; // @[Mux.scala 19:72:@26625.4]
  assign _T_30999 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,_T_30991}; // @[Mux.scala 19:72:@26626.4]
  assign _T_31001 = _T_2696 ? _T_30999 : 16'h0; // @[Mux.scala 19:72:@26627.4]
  assign _T_31016 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,_T_30879}; // @[Mux.scala 19:72:@26642.4]
  assign _T_31018 = _T_2697 ? _T_31016 : 16'h0; // @[Mux.scala 19:72:@26643.4]
  assign _T_31033 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,_T_30896}; // @[Mux.scala 19:72:@26658.4]
  assign _T_31035 = _T_2698 ? _T_31033 : 16'h0; // @[Mux.scala 19:72:@26659.4]
  assign _T_31050 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,_T_30913}; // @[Mux.scala 19:72:@26674.4]
  assign _T_31052 = _T_2699 ? _T_31050 : 16'h0; // @[Mux.scala 19:72:@26675.4]
  assign _T_31067 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,_T_30930}; // @[Mux.scala 19:72:@26690.4]
  assign _T_31069 = _T_2700 ? _T_31067 : 16'h0; // @[Mux.scala 19:72:@26691.4]
  assign _T_31084 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,_T_30947}; // @[Mux.scala 19:72:@26706.4]
  assign _T_31086 = _T_2701 ? _T_31084 : 16'h0; // @[Mux.scala 19:72:@26707.4]
  assign _T_31101 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,_T_30964}; // @[Mux.scala 19:72:@26722.4]
  assign _T_31103 = _T_2702 ? _T_31101 : 16'h0; // @[Mux.scala 19:72:@26723.4]
  assign _T_31118 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,_T_30981}; // @[Mux.scala 19:72:@26738.4]
  assign _T_31120 = _T_2703 ? _T_31118 : 16'h0; // @[Mux.scala 19:72:@26739.4]
  assign _T_31135 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,_T_30998}; // @[Mux.scala 19:72:@26754.4]
  assign _T_31137 = _T_2704 ? _T_31135 : 16'h0; // @[Mux.scala 19:72:@26755.4]
  assign _T_31138 = _T_30882 | _T_30899; // @[Mux.scala 19:72:@26756.4]
  assign _T_31139 = _T_31138 | _T_30916; // @[Mux.scala 19:72:@26757.4]
  assign _T_31140 = _T_31139 | _T_30933; // @[Mux.scala 19:72:@26758.4]
  assign _T_31141 = _T_31140 | _T_30950; // @[Mux.scala 19:72:@26759.4]
  assign _T_31142 = _T_31141 | _T_30967; // @[Mux.scala 19:72:@26760.4]
  assign _T_31143 = _T_31142 | _T_30984; // @[Mux.scala 19:72:@26761.4]
  assign _T_31144 = _T_31143 | _T_31001; // @[Mux.scala 19:72:@26762.4]
  assign _T_31145 = _T_31144 | _T_31018; // @[Mux.scala 19:72:@26763.4]
  assign _T_31146 = _T_31145 | _T_31035; // @[Mux.scala 19:72:@26764.4]
  assign _T_31147 = _T_31146 | _T_31052; // @[Mux.scala 19:72:@26765.4]
  assign _T_31148 = _T_31147 | _T_31069; // @[Mux.scala 19:72:@26766.4]
  assign _T_31149 = _T_31148 | _T_31086; // @[Mux.scala 19:72:@26767.4]
  assign _T_31150 = _T_31149 | _T_31103; // @[Mux.scala 19:72:@26768.4]
  assign _T_31151 = _T_31150 | _T_31120; // @[Mux.scala 19:72:@26769.4]
  assign _T_31152 = _T_31151 | _T_31137; // @[Mux.scala 19:72:@26770.4]
  assign _T_52326 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@27634.4]
  assign _T_52333 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8}; // @[Mux.scala 19:72:@27641.4]
  assign _T_52334 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,_T_52326}; // @[Mux.scala 19:72:@27642.4]
  assign _T_52336 = _T_2689 ? _T_52334 : 16'h0; // @[Mux.scala 19:72:@27643.4]
  assign _T_52343 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@27650.4]
  assign _T_52350 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9}; // @[Mux.scala 19:72:@27657.4]
  assign _T_52351 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,_T_52343}; // @[Mux.scala 19:72:@27658.4]
  assign _T_52353 = _T_2690 ? _T_52351 : 16'h0; // @[Mux.scala 19:72:@27659.4]
  assign _T_52360 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@27666.4]
  assign _T_52367 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10}; // @[Mux.scala 19:72:@27673.4]
  assign _T_52368 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,_T_52360}; // @[Mux.scala 19:72:@27674.4]
  assign _T_52370 = _T_2691 ? _T_52368 : 16'h0; // @[Mux.scala 19:72:@27675.4]
  assign _T_52377 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@27682.4]
  assign _T_52384 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11}; // @[Mux.scala 19:72:@27689.4]
  assign _T_52385 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,_T_52377}; // @[Mux.scala 19:72:@27690.4]
  assign _T_52387 = _T_2692 ? _T_52385 : 16'h0; // @[Mux.scala 19:72:@27691.4]
  assign _T_52394 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@27698.4]
  assign _T_52401 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12}; // @[Mux.scala 19:72:@27705.4]
  assign _T_52402 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,_T_52394}; // @[Mux.scala 19:72:@27706.4]
  assign _T_52404 = _T_2693 ? _T_52402 : 16'h0; // @[Mux.scala 19:72:@27707.4]
  assign _T_52411 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@27714.4]
  assign _T_52418 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13}; // @[Mux.scala 19:72:@27721.4]
  assign _T_52419 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,_T_52411}; // @[Mux.scala 19:72:@27722.4]
  assign _T_52421 = _T_2694 ? _T_52419 : 16'h0; // @[Mux.scala 19:72:@27723.4]
  assign _T_52428 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@27730.4]
  assign _T_52435 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14}; // @[Mux.scala 19:72:@27737.4]
  assign _T_52436 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,_T_52428}; // @[Mux.scala 19:72:@27738.4]
  assign _T_52438 = _T_2695 ? _T_52436 : 16'h0; // @[Mux.scala 19:72:@27739.4]
  assign _T_52445 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@27746.4]
  assign _T_52452 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15}; // @[Mux.scala 19:72:@27753.4]
  assign _T_52453 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,_T_52445}; // @[Mux.scala 19:72:@27754.4]
  assign _T_52455 = _T_2696 ? _T_52453 : 16'h0; // @[Mux.scala 19:72:@27755.4]
  assign _T_52470 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,_T_52333}; // @[Mux.scala 19:72:@27770.4]
  assign _T_52472 = _T_2697 ? _T_52470 : 16'h0; // @[Mux.scala 19:72:@27771.4]
  assign _T_52487 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,_T_52350}; // @[Mux.scala 19:72:@27786.4]
  assign _T_52489 = _T_2698 ? _T_52487 : 16'h0; // @[Mux.scala 19:72:@27787.4]
  assign _T_52504 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,_T_52367}; // @[Mux.scala 19:72:@27802.4]
  assign _T_52506 = _T_2699 ? _T_52504 : 16'h0; // @[Mux.scala 19:72:@27803.4]
  assign _T_52521 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,_T_52384}; // @[Mux.scala 19:72:@27818.4]
  assign _T_52523 = _T_2700 ? _T_52521 : 16'h0; // @[Mux.scala 19:72:@27819.4]
  assign _T_52538 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,_T_52401}; // @[Mux.scala 19:72:@27834.4]
  assign _T_52540 = _T_2701 ? _T_52538 : 16'h0; // @[Mux.scala 19:72:@27835.4]
  assign _T_52555 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,_T_52418}; // @[Mux.scala 19:72:@27850.4]
  assign _T_52557 = _T_2702 ? _T_52555 : 16'h0; // @[Mux.scala 19:72:@27851.4]
  assign _T_52572 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,_T_52435}; // @[Mux.scala 19:72:@27866.4]
  assign _T_52574 = _T_2703 ? _T_52572 : 16'h0; // @[Mux.scala 19:72:@27867.4]
  assign _T_52589 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,_T_52452}; // @[Mux.scala 19:72:@27882.4]
  assign _T_52591 = _T_2704 ? _T_52589 : 16'h0; // @[Mux.scala 19:72:@27883.4]
  assign _T_52592 = _T_52336 | _T_52353; // @[Mux.scala 19:72:@27884.4]
  assign _T_52593 = _T_52592 | _T_52370; // @[Mux.scala 19:72:@27885.4]
  assign _T_52594 = _T_52593 | _T_52387; // @[Mux.scala 19:72:@27886.4]
  assign _T_52595 = _T_52594 | _T_52404; // @[Mux.scala 19:72:@27887.4]
  assign _T_52596 = _T_52595 | _T_52421; // @[Mux.scala 19:72:@27888.4]
  assign _T_52597 = _T_52596 | _T_52438; // @[Mux.scala 19:72:@27889.4]
  assign _T_52598 = _T_52597 | _T_52455; // @[Mux.scala 19:72:@27890.4]
  assign _T_52599 = _T_52598 | _T_52472; // @[Mux.scala 19:72:@27891.4]
  assign _T_52600 = _T_52599 | _T_52489; // @[Mux.scala 19:72:@27892.4]
  assign _T_52601 = _T_52600 | _T_52506; // @[Mux.scala 19:72:@27893.4]
  assign _T_52602 = _T_52601 | _T_52523; // @[Mux.scala 19:72:@27894.4]
  assign _T_52603 = _T_52602 | _T_52540; // @[Mux.scala 19:72:@27895.4]
  assign _T_52604 = _T_52603 | _T_52557; // @[Mux.scala 19:72:@27896.4]
  assign _T_52605 = _T_52604 | _T_52574; // @[Mux.scala 19:72:@27897.4]
  assign _T_52606 = _T_52605 | _T_52591; // @[Mux.scala 19:72:@27898.4]
  assign _T_53184 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@28248.4]
  assign _T_53191 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8}; // @[Mux.scala 19:72:@28255.4]
  assign _T_53192 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,_T_53184}; // @[Mux.scala 19:72:@28256.4]
  assign _T_53194 = _T_2689 ? _T_53192 : 16'h0; // @[Mux.scala 19:72:@28257.4]
  assign _T_53201 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@28264.4]
  assign _T_53208 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9}; // @[Mux.scala 19:72:@28271.4]
  assign _T_53209 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,_T_53201}; // @[Mux.scala 19:72:@28272.4]
  assign _T_53211 = _T_2690 ? _T_53209 : 16'h0; // @[Mux.scala 19:72:@28273.4]
  assign _T_53218 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@28280.4]
  assign _T_53225 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10}; // @[Mux.scala 19:72:@28287.4]
  assign _T_53226 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,_T_53218}; // @[Mux.scala 19:72:@28288.4]
  assign _T_53228 = _T_2691 ? _T_53226 : 16'h0; // @[Mux.scala 19:72:@28289.4]
  assign _T_53235 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@28296.4]
  assign _T_53242 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11}; // @[Mux.scala 19:72:@28303.4]
  assign _T_53243 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,_T_53235}; // @[Mux.scala 19:72:@28304.4]
  assign _T_53245 = _T_2692 ? _T_53243 : 16'h0; // @[Mux.scala 19:72:@28305.4]
  assign _T_53252 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@28312.4]
  assign _T_53259 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12}; // @[Mux.scala 19:72:@28319.4]
  assign _T_53260 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,_T_53252}; // @[Mux.scala 19:72:@28320.4]
  assign _T_53262 = _T_2693 ? _T_53260 : 16'h0; // @[Mux.scala 19:72:@28321.4]
  assign _T_53269 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@28328.4]
  assign _T_53276 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13}; // @[Mux.scala 19:72:@28335.4]
  assign _T_53277 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,_T_53269}; // @[Mux.scala 19:72:@28336.4]
  assign _T_53279 = _T_2694 ? _T_53277 : 16'h0; // @[Mux.scala 19:72:@28337.4]
  assign _T_53286 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@28344.4]
  assign _T_53293 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14}; // @[Mux.scala 19:72:@28351.4]
  assign _T_53294 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,_T_53286}; // @[Mux.scala 19:72:@28352.4]
  assign _T_53296 = _T_2695 ? _T_53294 : 16'h0; // @[Mux.scala 19:72:@28353.4]
  assign _T_53303 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@28360.4]
  assign _T_53310 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15}; // @[Mux.scala 19:72:@28367.4]
  assign _T_53311 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,_T_53303}; // @[Mux.scala 19:72:@28368.4]
  assign _T_53313 = _T_2696 ? _T_53311 : 16'h0; // @[Mux.scala 19:72:@28369.4]
  assign _T_53328 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,_T_53191}; // @[Mux.scala 19:72:@28384.4]
  assign _T_53330 = _T_2697 ? _T_53328 : 16'h0; // @[Mux.scala 19:72:@28385.4]
  assign _T_53345 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,_T_53208}; // @[Mux.scala 19:72:@28400.4]
  assign _T_53347 = _T_2698 ? _T_53345 : 16'h0; // @[Mux.scala 19:72:@28401.4]
  assign _T_53362 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,_T_53225}; // @[Mux.scala 19:72:@28416.4]
  assign _T_53364 = _T_2699 ? _T_53362 : 16'h0; // @[Mux.scala 19:72:@28417.4]
  assign _T_53379 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,_T_53242}; // @[Mux.scala 19:72:@28432.4]
  assign _T_53381 = _T_2700 ? _T_53379 : 16'h0; // @[Mux.scala 19:72:@28433.4]
  assign _T_53396 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,_T_53259}; // @[Mux.scala 19:72:@28448.4]
  assign _T_53398 = _T_2701 ? _T_53396 : 16'h0; // @[Mux.scala 19:72:@28449.4]
  assign _T_53413 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,_T_53276}; // @[Mux.scala 19:72:@28464.4]
  assign _T_53415 = _T_2702 ? _T_53413 : 16'h0; // @[Mux.scala 19:72:@28465.4]
  assign _T_53430 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,_T_53293}; // @[Mux.scala 19:72:@28480.4]
  assign _T_53432 = _T_2703 ? _T_53430 : 16'h0; // @[Mux.scala 19:72:@28481.4]
  assign _T_53447 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,_T_53310}; // @[Mux.scala 19:72:@28496.4]
  assign _T_53449 = _T_2704 ? _T_53447 : 16'h0; // @[Mux.scala 19:72:@28497.4]
  assign _T_53450 = _T_53194 | _T_53211; // @[Mux.scala 19:72:@28498.4]
  assign _T_53451 = _T_53450 | _T_53228; // @[Mux.scala 19:72:@28499.4]
  assign _T_53452 = _T_53451 | _T_53245; // @[Mux.scala 19:72:@28500.4]
  assign _T_53453 = _T_53452 | _T_53262; // @[Mux.scala 19:72:@28501.4]
  assign _T_53454 = _T_53453 | _T_53279; // @[Mux.scala 19:72:@28502.4]
  assign _T_53455 = _T_53454 | _T_53296; // @[Mux.scala 19:72:@28503.4]
  assign _T_53456 = _T_53455 | _T_53313; // @[Mux.scala 19:72:@28504.4]
  assign _T_53457 = _T_53456 | _T_53330; // @[Mux.scala 19:72:@28505.4]
  assign _T_53458 = _T_53457 | _T_53347; // @[Mux.scala 19:72:@28506.4]
  assign _T_53459 = _T_53458 | _T_53364; // @[Mux.scala 19:72:@28507.4]
  assign _T_53460 = _T_53459 | _T_53381; // @[Mux.scala 19:72:@28508.4]
  assign _T_53461 = _T_53460 | _T_53398; // @[Mux.scala 19:72:@28509.4]
  assign _T_53462 = _T_53461 | _T_53415; // @[Mux.scala 19:72:@28510.4]
  assign _T_53463 = _T_53462 | _T_53432; // @[Mux.scala 19:72:@28511.4]
  assign _T_53464 = _T_53463 | _T_53449; // @[Mux.scala 19:72:@28512.4]
  assign _T_54042 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@28862.4]
  assign _T_54049 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8}; // @[Mux.scala 19:72:@28869.4]
  assign _T_54050 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,_T_54042}; // @[Mux.scala 19:72:@28870.4]
  assign _T_54052 = _T_2689 ? _T_54050 : 16'h0; // @[Mux.scala 19:72:@28871.4]
  assign _T_54059 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@28878.4]
  assign _T_54066 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9}; // @[Mux.scala 19:72:@28885.4]
  assign _T_54067 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,_T_54059}; // @[Mux.scala 19:72:@28886.4]
  assign _T_54069 = _T_2690 ? _T_54067 : 16'h0; // @[Mux.scala 19:72:@28887.4]
  assign _T_54076 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@28894.4]
  assign _T_54083 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10}; // @[Mux.scala 19:72:@28901.4]
  assign _T_54084 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,_T_54076}; // @[Mux.scala 19:72:@28902.4]
  assign _T_54086 = _T_2691 ? _T_54084 : 16'h0; // @[Mux.scala 19:72:@28903.4]
  assign _T_54093 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@28910.4]
  assign _T_54100 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11}; // @[Mux.scala 19:72:@28917.4]
  assign _T_54101 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,_T_54093}; // @[Mux.scala 19:72:@28918.4]
  assign _T_54103 = _T_2692 ? _T_54101 : 16'h0; // @[Mux.scala 19:72:@28919.4]
  assign _T_54110 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@28926.4]
  assign _T_54117 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12}; // @[Mux.scala 19:72:@28933.4]
  assign _T_54118 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,_T_54110}; // @[Mux.scala 19:72:@28934.4]
  assign _T_54120 = _T_2693 ? _T_54118 : 16'h0; // @[Mux.scala 19:72:@28935.4]
  assign _T_54127 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@28942.4]
  assign _T_54134 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13}; // @[Mux.scala 19:72:@28949.4]
  assign _T_54135 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,_T_54127}; // @[Mux.scala 19:72:@28950.4]
  assign _T_54137 = _T_2694 ? _T_54135 : 16'h0; // @[Mux.scala 19:72:@28951.4]
  assign _T_54144 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@28958.4]
  assign _T_54151 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14}; // @[Mux.scala 19:72:@28965.4]
  assign _T_54152 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,_T_54144}; // @[Mux.scala 19:72:@28966.4]
  assign _T_54154 = _T_2695 ? _T_54152 : 16'h0; // @[Mux.scala 19:72:@28967.4]
  assign _T_54161 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@28974.4]
  assign _T_54168 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15}; // @[Mux.scala 19:72:@28981.4]
  assign _T_54169 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,_T_54161}; // @[Mux.scala 19:72:@28982.4]
  assign _T_54171 = _T_2696 ? _T_54169 : 16'h0; // @[Mux.scala 19:72:@28983.4]
  assign _T_54186 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,_T_54049}; // @[Mux.scala 19:72:@28998.4]
  assign _T_54188 = _T_2697 ? _T_54186 : 16'h0; // @[Mux.scala 19:72:@28999.4]
  assign _T_54203 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,_T_54066}; // @[Mux.scala 19:72:@29014.4]
  assign _T_54205 = _T_2698 ? _T_54203 : 16'h0; // @[Mux.scala 19:72:@29015.4]
  assign _T_54220 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,_T_54083}; // @[Mux.scala 19:72:@29030.4]
  assign _T_54222 = _T_2699 ? _T_54220 : 16'h0; // @[Mux.scala 19:72:@29031.4]
  assign _T_54237 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,_T_54100}; // @[Mux.scala 19:72:@29046.4]
  assign _T_54239 = _T_2700 ? _T_54237 : 16'h0; // @[Mux.scala 19:72:@29047.4]
  assign _T_54254 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,_T_54117}; // @[Mux.scala 19:72:@29062.4]
  assign _T_54256 = _T_2701 ? _T_54254 : 16'h0; // @[Mux.scala 19:72:@29063.4]
  assign _T_54271 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,_T_54134}; // @[Mux.scala 19:72:@29078.4]
  assign _T_54273 = _T_2702 ? _T_54271 : 16'h0; // @[Mux.scala 19:72:@29079.4]
  assign _T_54288 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,_T_54151}; // @[Mux.scala 19:72:@29094.4]
  assign _T_54290 = _T_2703 ? _T_54288 : 16'h0; // @[Mux.scala 19:72:@29095.4]
  assign _T_54305 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,_T_54168}; // @[Mux.scala 19:72:@29110.4]
  assign _T_54307 = _T_2704 ? _T_54305 : 16'h0; // @[Mux.scala 19:72:@29111.4]
  assign _T_54308 = _T_54052 | _T_54069; // @[Mux.scala 19:72:@29112.4]
  assign _T_54309 = _T_54308 | _T_54086; // @[Mux.scala 19:72:@29113.4]
  assign _T_54310 = _T_54309 | _T_54103; // @[Mux.scala 19:72:@29114.4]
  assign _T_54311 = _T_54310 | _T_54120; // @[Mux.scala 19:72:@29115.4]
  assign _T_54312 = _T_54311 | _T_54137; // @[Mux.scala 19:72:@29116.4]
  assign _T_54313 = _T_54312 | _T_54154; // @[Mux.scala 19:72:@29117.4]
  assign _T_54314 = _T_54313 | _T_54171; // @[Mux.scala 19:72:@29118.4]
  assign _T_54315 = _T_54314 | _T_54188; // @[Mux.scala 19:72:@29119.4]
  assign _T_54316 = _T_54315 | _T_54205; // @[Mux.scala 19:72:@29120.4]
  assign _T_54317 = _T_54316 | _T_54222; // @[Mux.scala 19:72:@29121.4]
  assign _T_54318 = _T_54317 | _T_54239; // @[Mux.scala 19:72:@29122.4]
  assign _T_54319 = _T_54318 | _T_54256; // @[Mux.scala 19:72:@29123.4]
  assign _T_54320 = _T_54319 | _T_54273; // @[Mux.scala 19:72:@29124.4]
  assign _T_54321 = _T_54320 | _T_54290; // @[Mux.scala 19:72:@29125.4]
  assign _T_54322 = _T_54321 | _T_54307; // @[Mux.scala 19:72:@29126.4]
  assign _T_54900 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@29476.4]
  assign _T_54907 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8}; // @[Mux.scala 19:72:@29483.4]
  assign _T_54908 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,_T_54900}; // @[Mux.scala 19:72:@29484.4]
  assign _T_54910 = _T_2689 ? _T_54908 : 16'h0; // @[Mux.scala 19:72:@29485.4]
  assign _T_54917 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@29492.4]
  assign _T_54924 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9}; // @[Mux.scala 19:72:@29499.4]
  assign _T_54925 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,_T_54917}; // @[Mux.scala 19:72:@29500.4]
  assign _T_54927 = _T_2690 ? _T_54925 : 16'h0; // @[Mux.scala 19:72:@29501.4]
  assign _T_54934 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@29508.4]
  assign _T_54941 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10}; // @[Mux.scala 19:72:@29515.4]
  assign _T_54942 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,_T_54934}; // @[Mux.scala 19:72:@29516.4]
  assign _T_54944 = _T_2691 ? _T_54942 : 16'h0; // @[Mux.scala 19:72:@29517.4]
  assign _T_54951 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@29524.4]
  assign _T_54958 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11}; // @[Mux.scala 19:72:@29531.4]
  assign _T_54959 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,_T_54951}; // @[Mux.scala 19:72:@29532.4]
  assign _T_54961 = _T_2692 ? _T_54959 : 16'h0; // @[Mux.scala 19:72:@29533.4]
  assign _T_54968 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@29540.4]
  assign _T_54975 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12}; // @[Mux.scala 19:72:@29547.4]
  assign _T_54976 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,_T_54968}; // @[Mux.scala 19:72:@29548.4]
  assign _T_54978 = _T_2693 ? _T_54976 : 16'h0; // @[Mux.scala 19:72:@29549.4]
  assign _T_54985 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@29556.4]
  assign _T_54992 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13}; // @[Mux.scala 19:72:@29563.4]
  assign _T_54993 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,_T_54985}; // @[Mux.scala 19:72:@29564.4]
  assign _T_54995 = _T_2694 ? _T_54993 : 16'h0; // @[Mux.scala 19:72:@29565.4]
  assign _T_55002 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@29572.4]
  assign _T_55009 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14}; // @[Mux.scala 19:72:@29579.4]
  assign _T_55010 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,_T_55002}; // @[Mux.scala 19:72:@29580.4]
  assign _T_55012 = _T_2695 ? _T_55010 : 16'h0; // @[Mux.scala 19:72:@29581.4]
  assign _T_55019 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@29588.4]
  assign _T_55026 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15}; // @[Mux.scala 19:72:@29595.4]
  assign _T_55027 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,_T_55019}; // @[Mux.scala 19:72:@29596.4]
  assign _T_55029 = _T_2696 ? _T_55027 : 16'h0; // @[Mux.scala 19:72:@29597.4]
  assign _T_55044 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,_T_54907}; // @[Mux.scala 19:72:@29612.4]
  assign _T_55046 = _T_2697 ? _T_55044 : 16'h0; // @[Mux.scala 19:72:@29613.4]
  assign _T_55061 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,_T_54924}; // @[Mux.scala 19:72:@29628.4]
  assign _T_55063 = _T_2698 ? _T_55061 : 16'h0; // @[Mux.scala 19:72:@29629.4]
  assign _T_55078 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,_T_54941}; // @[Mux.scala 19:72:@29644.4]
  assign _T_55080 = _T_2699 ? _T_55078 : 16'h0; // @[Mux.scala 19:72:@29645.4]
  assign _T_55095 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,_T_54958}; // @[Mux.scala 19:72:@29660.4]
  assign _T_55097 = _T_2700 ? _T_55095 : 16'h0; // @[Mux.scala 19:72:@29661.4]
  assign _T_55112 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,_T_54975}; // @[Mux.scala 19:72:@29676.4]
  assign _T_55114 = _T_2701 ? _T_55112 : 16'h0; // @[Mux.scala 19:72:@29677.4]
  assign _T_55129 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,_T_54992}; // @[Mux.scala 19:72:@29692.4]
  assign _T_55131 = _T_2702 ? _T_55129 : 16'h0; // @[Mux.scala 19:72:@29693.4]
  assign _T_55146 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,_T_55009}; // @[Mux.scala 19:72:@29708.4]
  assign _T_55148 = _T_2703 ? _T_55146 : 16'h0; // @[Mux.scala 19:72:@29709.4]
  assign _T_55163 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,_T_55026}; // @[Mux.scala 19:72:@29724.4]
  assign _T_55165 = _T_2704 ? _T_55163 : 16'h0; // @[Mux.scala 19:72:@29725.4]
  assign _T_55166 = _T_54910 | _T_54927; // @[Mux.scala 19:72:@29726.4]
  assign _T_55167 = _T_55166 | _T_54944; // @[Mux.scala 19:72:@29727.4]
  assign _T_55168 = _T_55167 | _T_54961; // @[Mux.scala 19:72:@29728.4]
  assign _T_55169 = _T_55168 | _T_54978; // @[Mux.scala 19:72:@29729.4]
  assign _T_55170 = _T_55169 | _T_54995; // @[Mux.scala 19:72:@29730.4]
  assign _T_55171 = _T_55170 | _T_55012; // @[Mux.scala 19:72:@29731.4]
  assign _T_55172 = _T_55171 | _T_55029; // @[Mux.scala 19:72:@29732.4]
  assign _T_55173 = _T_55172 | _T_55046; // @[Mux.scala 19:72:@29733.4]
  assign _T_55174 = _T_55173 | _T_55063; // @[Mux.scala 19:72:@29734.4]
  assign _T_55175 = _T_55174 | _T_55080; // @[Mux.scala 19:72:@29735.4]
  assign _T_55176 = _T_55175 | _T_55097; // @[Mux.scala 19:72:@29736.4]
  assign _T_55177 = _T_55176 | _T_55114; // @[Mux.scala 19:72:@29737.4]
  assign _T_55178 = _T_55177 | _T_55131; // @[Mux.scala 19:72:@29738.4]
  assign _T_55179 = _T_55178 | _T_55148; // @[Mux.scala 19:72:@29739.4]
  assign _T_55180 = _T_55179 | _T_55165; // @[Mux.scala 19:72:@29740.4]
  assign _T_55758 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@30090.4]
  assign _T_55765 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8}; // @[Mux.scala 19:72:@30097.4]
  assign _T_55766 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,_T_55758}; // @[Mux.scala 19:72:@30098.4]
  assign _T_55768 = _T_2689 ? _T_55766 : 16'h0; // @[Mux.scala 19:72:@30099.4]
  assign _T_55775 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@30106.4]
  assign _T_55782 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9}; // @[Mux.scala 19:72:@30113.4]
  assign _T_55783 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,_T_55775}; // @[Mux.scala 19:72:@30114.4]
  assign _T_55785 = _T_2690 ? _T_55783 : 16'h0; // @[Mux.scala 19:72:@30115.4]
  assign _T_55792 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@30122.4]
  assign _T_55799 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10}; // @[Mux.scala 19:72:@30129.4]
  assign _T_55800 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,_T_55792}; // @[Mux.scala 19:72:@30130.4]
  assign _T_55802 = _T_2691 ? _T_55800 : 16'h0; // @[Mux.scala 19:72:@30131.4]
  assign _T_55809 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@30138.4]
  assign _T_55816 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11}; // @[Mux.scala 19:72:@30145.4]
  assign _T_55817 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,_T_55809}; // @[Mux.scala 19:72:@30146.4]
  assign _T_55819 = _T_2692 ? _T_55817 : 16'h0; // @[Mux.scala 19:72:@30147.4]
  assign _T_55826 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@30154.4]
  assign _T_55833 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12}; // @[Mux.scala 19:72:@30161.4]
  assign _T_55834 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,_T_55826}; // @[Mux.scala 19:72:@30162.4]
  assign _T_55836 = _T_2693 ? _T_55834 : 16'h0; // @[Mux.scala 19:72:@30163.4]
  assign _T_55843 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@30170.4]
  assign _T_55850 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13}; // @[Mux.scala 19:72:@30177.4]
  assign _T_55851 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,_T_55843}; // @[Mux.scala 19:72:@30178.4]
  assign _T_55853 = _T_2694 ? _T_55851 : 16'h0; // @[Mux.scala 19:72:@30179.4]
  assign _T_55860 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@30186.4]
  assign _T_55867 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14}; // @[Mux.scala 19:72:@30193.4]
  assign _T_55868 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,_T_55860}; // @[Mux.scala 19:72:@30194.4]
  assign _T_55870 = _T_2695 ? _T_55868 : 16'h0; // @[Mux.scala 19:72:@30195.4]
  assign _T_55877 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@30202.4]
  assign _T_55884 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15}; // @[Mux.scala 19:72:@30209.4]
  assign _T_55885 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,_T_55877}; // @[Mux.scala 19:72:@30210.4]
  assign _T_55887 = _T_2696 ? _T_55885 : 16'h0; // @[Mux.scala 19:72:@30211.4]
  assign _T_55902 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,_T_55765}; // @[Mux.scala 19:72:@30226.4]
  assign _T_55904 = _T_2697 ? _T_55902 : 16'h0; // @[Mux.scala 19:72:@30227.4]
  assign _T_55919 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,_T_55782}; // @[Mux.scala 19:72:@30242.4]
  assign _T_55921 = _T_2698 ? _T_55919 : 16'h0; // @[Mux.scala 19:72:@30243.4]
  assign _T_55936 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,_T_55799}; // @[Mux.scala 19:72:@30258.4]
  assign _T_55938 = _T_2699 ? _T_55936 : 16'h0; // @[Mux.scala 19:72:@30259.4]
  assign _T_55953 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,_T_55816}; // @[Mux.scala 19:72:@30274.4]
  assign _T_55955 = _T_2700 ? _T_55953 : 16'h0; // @[Mux.scala 19:72:@30275.4]
  assign _T_55970 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,_T_55833}; // @[Mux.scala 19:72:@30290.4]
  assign _T_55972 = _T_2701 ? _T_55970 : 16'h0; // @[Mux.scala 19:72:@30291.4]
  assign _T_55987 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,_T_55850}; // @[Mux.scala 19:72:@30306.4]
  assign _T_55989 = _T_2702 ? _T_55987 : 16'h0; // @[Mux.scala 19:72:@30307.4]
  assign _T_56004 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,_T_55867}; // @[Mux.scala 19:72:@30322.4]
  assign _T_56006 = _T_2703 ? _T_56004 : 16'h0; // @[Mux.scala 19:72:@30323.4]
  assign _T_56021 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,_T_55884}; // @[Mux.scala 19:72:@30338.4]
  assign _T_56023 = _T_2704 ? _T_56021 : 16'h0; // @[Mux.scala 19:72:@30339.4]
  assign _T_56024 = _T_55768 | _T_55785; // @[Mux.scala 19:72:@30340.4]
  assign _T_56025 = _T_56024 | _T_55802; // @[Mux.scala 19:72:@30341.4]
  assign _T_56026 = _T_56025 | _T_55819; // @[Mux.scala 19:72:@30342.4]
  assign _T_56027 = _T_56026 | _T_55836; // @[Mux.scala 19:72:@30343.4]
  assign _T_56028 = _T_56027 | _T_55853; // @[Mux.scala 19:72:@30344.4]
  assign _T_56029 = _T_56028 | _T_55870; // @[Mux.scala 19:72:@30345.4]
  assign _T_56030 = _T_56029 | _T_55887; // @[Mux.scala 19:72:@30346.4]
  assign _T_56031 = _T_56030 | _T_55904; // @[Mux.scala 19:72:@30347.4]
  assign _T_56032 = _T_56031 | _T_55921; // @[Mux.scala 19:72:@30348.4]
  assign _T_56033 = _T_56032 | _T_55938; // @[Mux.scala 19:72:@30349.4]
  assign _T_56034 = _T_56033 | _T_55955; // @[Mux.scala 19:72:@30350.4]
  assign _T_56035 = _T_56034 | _T_55972; // @[Mux.scala 19:72:@30351.4]
  assign _T_56036 = _T_56035 | _T_55989; // @[Mux.scala 19:72:@30352.4]
  assign _T_56037 = _T_56036 | _T_56006; // @[Mux.scala 19:72:@30353.4]
  assign _T_56038 = _T_56037 | _T_56023; // @[Mux.scala 19:72:@30354.4]
  assign _T_56616 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@30704.4]
  assign _T_56623 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8}; // @[Mux.scala 19:72:@30711.4]
  assign _T_56624 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,_T_56616}; // @[Mux.scala 19:72:@30712.4]
  assign _T_56626 = _T_2689 ? _T_56624 : 16'h0; // @[Mux.scala 19:72:@30713.4]
  assign _T_56633 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@30720.4]
  assign _T_56640 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9}; // @[Mux.scala 19:72:@30727.4]
  assign _T_56641 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,_T_56633}; // @[Mux.scala 19:72:@30728.4]
  assign _T_56643 = _T_2690 ? _T_56641 : 16'h0; // @[Mux.scala 19:72:@30729.4]
  assign _T_56650 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@30736.4]
  assign _T_56657 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10}; // @[Mux.scala 19:72:@30743.4]
  assign _T_56658 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,_T_56650}; // @[Mux.scala 19:72:@30744.4]
  assign _T_56660 = _T_2691 ? _T_56658 : 16'h0; // @[Mux.scala 19:72:@30745.4]
  assign _T_56667 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@30752.4]
  assign _T_56674 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11}; // @[Mux.scala 19:72:@30759.4]
  assign _T_56675 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,_T_56667}; // @[Mux.scala 19:72:@30760.4]
  assign _T_56677 = _T_2692 ? _T_56675 : 16'h0; // @[Mux.scala 19:72:@30761.4]
  assign _T_56684 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@30768.4]
  assign _T_56691 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12}; // @[Mux.scala 19:72:@30775.4]
  assign _T_56692 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,_T_56684}; // @[Mux.scala 19:72:@30776.4]
  assign _T_56694 = _T_2693 ? _T_56692 : 16'h0; // @[Mux.scala 19:72:@30777.4]
  assign _T_56701 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@30784.4]
  assign _T_56708 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13}; // @[Mux.scala 19:72:@30791.4]
  assign _T_56709 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,_T_56701}; // @[Mux.scala 19:72:@30792.4]
  assign _T_56711 = _T_2694 ? _T_56709 : 16'h0; // @[Mux.scala 19:72:@30793.4]
  assign _T_56718 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@30800.4]
  assign _T_56725 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14}; // @[Mux.scala 19:72:@30807.4]
  assign _T_56726 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,_T_56718}; // @[Mux.scala 19:72:@30808.4]
  assign _T_56728 = _T_2695 ? _T_56726 : 16'h0; // @[Mux.scala 19:72:@30809.4]
  assign _T_56735 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@30816.4]
  assign _T_56742 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15}; // @[Mux.scala 19:72:@30823.4]
  assign _T_56743 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,_T_56735}; // @[Mux.scala 19:72:@30824.4]
  assign _T_56745 = _T_2696 ? _T_56743 : 16'h0; // @[Mux.scala 19:72:@30825.4]
  assign _T_56760 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,_T_56623}; // @[Mux.scala 19:72:@30840.4]
  assign _T_56762 = _T_2697 ? _T_56760 : 16'h0; // @[Mux.scala 19:72:@30841.4]
  assign _T_56777 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,_T_56640}; // @[Mux.scala 19:72:@30856.4]
  assign _T_56779 = _T_2698 ? _T_56777 : 16'h0; // @[Mux.scala 19:72:@30857.4]
  assign _T_56794 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,_T_56657}; // @[Mux.scala 19:72:@30872.4]
  assign _T_56796 = _T_2699 ? _T_56794 : 16'h0; // @[Mux.scala 19:72:@30873.4]
  assign _T_56811 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,_T_56674}; // @[Mux.scala 19:72:@30888.4]
  assign _T_56813 = _T_2700 ? _T_56811 : 16'h0; // @[Mux.scala 19:72:@30889.4]
  assign _T_56828 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,_T_56691}; // @[Mux.scala 19:72:@30904.4]
  assign _T_56830 = _T_2701 ? _T_56828 : 16'h0; // @[Mux.scala 19:72:@30905.4]
  assign _T_56845 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,_T_56708}; // @[Mux.scala 19:72:@30920.4]
  assign _T_56847 = _T_2702 ? _T_56845 : 16'h0; // @[Mux.scala 19:72:@30921.4]
  assign _T_56862 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,_T_56725}; // @[Mux.scala 19:72:@30936.4]
  assign _T_56864 = _T_2703 ? _T_56862 : 16'h0; // @[Mux.scala 19:72:@30937.4]
  assign _T_56879 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,_T_56742}; // @[Mux.scala 19:72:@30952.4]
  assign _T_56881 = _T_2704 ? _T_56879 : 16'h0; // @[Mux.scala 19:72:@30953.4]
  assign _T_56882 = _T_56626 | _T_56643; // @[Mux.scala 19:72:@30954.4]
  assign _T_56883 = _T_56882 | _T_56660; // @[Mux.scala 19:72:@30955.4]
  assign _T_56884 = _T_56883 | _T_56677; // @[Mux.scala 19:72:@30956.4]
  assign _T_56885 = _T_56884 | _T_56694; // @[Mux.scala 19:72:@30957.4]
  assign _T_56886 = _T_56885 | _T_56711; // @[Mux.scala 19:72:@30958.4]
  assign _T_56887 = _T_56886 | _T_56728; // @[Mux.scala 19:72:@30959.4]
  assign _T_56888 = _T_56887 | _T_56745; // @[Mux.scala 19:72:@30960.4]
  assign _T_56889 = _T_56888 | _T_56762; // @[Mux.scala 19:72:@30961.4]
  assign _T_56890 = _T_56889 | _T_56779; // @[Mux.scala 19:72:@30962.4]
  assign _T_56891 = _T_56890 | _T_56796; // @[Mux.scala 19:72:@30963.4]
  assign _T_56892 = _T_56891 | _T_56813; // @[Mux.scala 19:72:@30964.4]
  assign _T_56893 = _T_56892 | _T_56830; // @[Mux.scala 19:72:@30965.4]
  assign _T_56894 = _T_56893 | _T_56847; // @[Mux.scala 19:72:@30966.4]
  assign _T_56895 = _T_56894 | _T_56864; // @[Mux.scala 19:72:@30967.4]
  assign _T_56896 = _T_56895 | _T_56881; // @[Mux.scala 19:72:@30968.4]
  assign _T_57474 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@31318.4]
  assign _T_57481 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8}; // @[Mux.scala 19:72:@31325.4]
  assign _T_57482 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,_T_57474}; // @[Mux.scala 19:72:@31326.4]
  assign _T_57484 = _T_2689 ? _T_57482 : 16'h0; // @[Mux.scala 19:72:@31327.4]
  assign _T_57491 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@31334.4]
  assign _T_57498 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9}; // @[Mux.scala 19:72:@31341.4]
  assign _T_57499 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,_T_57491}; // @[Mux.scala 19:72:@31342.4]
  assign _T_57501 = _T_2690 ? _T_57499 : 16'h0; // @[Mux.scala 19:72:@31343.4]
  assign _T_57508 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@31350.4]
  assign _T_57515 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10}; // @[Mux.scala 19:72:@31357.4]
  assign _T_57516 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,_T_57508}; // @[Mux.scala 19:72:@31358.4]
  assign _T_57518 = _T_2691 ? _T_57516 : 16'h0; // @[Mux.scala 19:72:@31359.4]
  assign _T_57525 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@31366.4]
  assign _T_57532 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11}; // @[Mux.scala 19:72:@31373.4]
  assign _T_57533 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,_T_57525}; // @[Mux.scala 19:72:@31374.4]
  assign _T_57535 = _T_2692 ? _T_57533 : 16'h0; // @[Mux.scala 19:72:@31375.4]
  assign _T_57542 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@31382.4]
  assign _T_57549 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12}; // @[Mux.scala 19:72:@31389.4]
  assign _T_57550 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,_T_57542}; // @[Mux.scala 19:72:@31390.4]
  assign _T_57552 = _T_2693 ? _T_57550 : 16'h0; // @[Mux.scala 19:72:@31391.4]
  assign _T_57559 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@31398.4]
  assign _T_57566 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13}; // @[Mux.scala 19:72:@31405.4]
  assign _T_57567 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,_T_57559}; // @[Mux.scala 19:72:@31406.4]
  assign _T_57569 = _T_2694 ? _T_57567 : 16'h0; // @[Mux.scala 19:72:@31407.4]
  assign _T_57576 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@31414.4]
  assign _T_57583 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14}; // @[Mux.scala 19:72:@31421.4]
  assign _T_57584 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,_T_57576}; // @[Mux.scala 19:72:@31422.4]
  assign _T_57586 = _T_2695 ? _T_57584 : 16'h0; // @[Mux.scala 19:72:@31423.4]
  assign _T_57593 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@31430.4]
  assign _T_57600 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15}; // @[Mux.scala 19:72:@31437.4]
  assign _T_57601 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,_T_57593}; // @[Mux.scala 19:72:@31438.4]
  assign _T_57603 = _T_2696 ? _T_57601 : 16'h0; // @[Mux.scala 19:72:@31439.4]
  assign _T_57618 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,_T_57481}; // @[Mux.scala 19:72:@31454.4]
  assign _T_57620 = _T_2697 ? _T_57618 : 16'h0; // @[Mux.scala 19:72:@31455.4]
  assign _T_57635 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,_T_57498}; // @[Mux.scala 19:72:@31470.4]
  assign _T_57637 = _T_2698 ? _T_57635 : 16'h0; // @[Mux.scala 19:72:@31471.4]
  assign _T_57652 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,_T_57515}; // @[Mux.scala 19:72:@31486.4]
  assign _T_57654 = _T_2699 ? _T_57652 : 16'h0; // @[Mux.scala 19:72:@31487.4]
  assign _T_57669 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,_T_57532}; // @[Mux.scala 19:72:@31502.4]
  assign _T_57671 = _T_2700 ? _T_57669 : 16'h0; // @[Mux.scala 19:72:@31503.4]
  assign _T_57686 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,_T_57549}; // @[Mux.scala 19:72:@31518.4]
  assign _T_57688 = _T_2701 ? _T_57686 : 16'h0; // @[Mux.scala 19:72:@31519.4]
  assign _T_57703 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,_T_57566}; // @[Mux.scala 19:72:@31534.4]
  assign _T_57705 = _T_2702 ? _T_57703 : 16'h0; // @[Mux.scala 19:72:@31535.4]
  assign _T_57720 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,_T_57583}; // @[Mux.scala 19:72:@31550.4]
  assign _T_57722 = _T_2703 ? _T_57720 : 16'h0; // @[Mux.scala 19:72:@31551.4]
  assign _T_57737 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,_T_57600}; // @[Mux.scala 19:72:@31566.4]
  assign _T_57739 = _T_2704 ? _T_57737 : 16'h0; // @[Mux.scala 19:72:@31567.4]
  assign _T_57740 = _T_57484 | _T_57501; // @[Mux.scala 19:72:@31568.4]
  assign _T_57741 = _T_57740 | _T_57518; // @[Mux.scala 19:72:@31569.4]
  assign _T_57742 = _T_57741 | _T_57535; // @[Mux.scala 19:72:@31570.4]
  assign _T_57743 = _T_57742 | _T_57552; // @[Mux.scala 19:72:@31571.4]
  assign _T_57744 = _T_57743 | _T_57569; // @[Mux.scala 19:72:@31572.4]
  assign _T_57745 = _T_57744 | _T_57586; // @[Mux.scala 19:72:@31573.4]
  assign _T_57746 = _T_57745 | _T_57603; // @[Mux.scala 19:72:@31574.4]
  assign _T_57747 = _T_57746 | _T_57620; // @[Mux.scala 19:72:@31575.4]
  assign _T_57748 = _T_57747 | _T_57637; // @[Mux.scala 19:72:@31576.4]
  assign _T_57749 = _T_57748 | _T_57654; // @[Mux.scala 19:72:@31577.4]
  assign _T_57750 = _T_57749 | _T_57671; // @[Mux.scala 19:72:@31578.4]
  assign _T_57751 = _T_57750 | _T_57688; // @[Mux.scala 19:72:@31579.4]
  assign _T_57752 = _T_57751 | _T_57705; // @[Mux.scala 19:72:@31580.4]
  assign _T_57753 = _T_57752 | _T_57722; // @[Mux.scala 19:72:@31581.4]
  assign _T_57754 = _T_57753 | _T_57739; // @[Mux.scala 19:72:@31582.4]
  assign _T_58332 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@31932.4]
  assign _T_58339 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8}; // @[Mux.scala 19:72:@31939.4]
  assign _T_58340 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,_T_58332}; // @[Mux.scala 19:72:@31940.4]
  assign _T_58342 = _T_2689 ? _T_58340 : 16'h0; // @[Mux.scala 19:72:@31941.4]
  assign _T_58349 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@31948.4]
  assign _T_58356 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9}; // @[Mux.scala 19:72:@31955.4]
  assign _T_58357 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,_T_58349}; // @[Mux.scala 19:72:@31956.4]
  assign _T_58359 = _T_2690 ? _T_58357 : 16'h0; // @[Mux.scala 19:72:@31957.4]
  assign _T_58366 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@31964.4]
  assign _T_58373 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10}; // @[Mux.scala 19:72:@31971.4]
  assign _T_58374 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,_T_58366}; // @[Mux.scala 19:72:@31972.4]
  assign _T_58376 = _T_2691 ? _T_58374 : 16'h0; // @[Mux.scala 19:72:@31973.4]
  assign _T_58383 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@31980.4]
  assign _T_58390 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11}; // @[Mux.scala 19:72:@31987.4]
  assign _T_58391 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,_T_58383}; // @[Mux.scala 19:72:@31988.4]
  assign _T_58393 = _T_2692 ? _T_58391 : 16'h0; // @[Mux.scala 19:72:@31989.4]
  assign _T_58400 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@31996.4]
  assign _T_58407 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12}; // @[Mux.scala 19:72:@32003.4]
  assign _T_58408 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,_T_58400}; // @[Mux.scala 19:72:@32004.4]
  assign _T_58410 = _T_2693 ? _T_58408 : 16'h0; // @[Mux.scala 19:72:@32005.4]
  assign _T_58417 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@32012.4]
  assign _T_58424 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13}; // @[Mux.scala 19:72:@32019.4]
  assign _T_58425 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,_T_58417}; // @[Mux.scala 19:72:@32020.4]
  assign _T_58427 = _T_2694 ? _T_58425 : 16'h0; // @[Mux.scala 19:72:@32021.4]
  assign _T_58434 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@32028.4]
  assign _T_58441 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14}; // @[Mux.scala 19:72:@32035.4]
  assign _T_58442 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,_T_58434}; // @[Mux.scala 19:72:@32036.4]
  assign _T_58444 = _T_2695 ? _T_58442 : 16'h0; // @[Mux.scala 19:72:@32037.4]
  assign _T_58451 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@32044.4]
  assign _T_58458 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15}; // @[Mux.scala 19:72:@32051.4]
  assign _T_58459 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,_T_58451}; // @[Mux.scala 19:72:@32052.4]
  assign _T_58461 = _T_2696 ? _T_58459 : 16'h0; // @[Mux.scala 19:72:@32053.4]
  assign _T_58476 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,_T_58339}; // @[Mux.scala 19:72:@32068.4]
  assign _T_58478 = _T_2697 ? _T_58476 : 16'h0; // @[Mux.scala 19:72:@32069.4]
  assign _T_58493 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,_T_58356}; // @[Mux.scala 19:72:@32084.4]
  assign _T_58495 = _T_2698 ? _T_58493 : 16'h0; // @[Mux.scala 19:72:@32085.4]
  assign _T_58510 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,_T_58373}; // @[Mux.scala 19:72:@32100.4]
  assign _T_58512 = _T_2699 ? _T_58510 : 16'h0; // @[Mux.scala 19:72:@32101.4]
  assign _T_58527 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,_T_58390}; // @[Mux.scala 19:72:@32116.4]
  assign _T_58529 = _T_2700 ? _T_58527 : 16'h0; // @[Mux.scala 19:72:@32117.4]
  assign _T_58544 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,_T_58407}; // @[Mux.scala 19:72:@32132.4]
  assign _T_58546 = _T_2701 ? _T_58544 : 16'h0; // @[Mux.scala 19:72:@32133.4]
  assign _T_58561 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,_T_58424}; // @[Mux.scala 19:72:@32148.4]
  assign _T_58563 = _T_2702 ? _T_58561 : 16'h0; // @[Mux.scala 19:72:@32149.4]
  assign _T_58578 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,_T_58441}; // @[Mux.scala 19:72:@32164.4]
  assign _T_58580 = _T_2703 ? _T_58578 : 16'h0; // @[Mux.scala 19:72:@32165.4]
  assign _T_58595 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,_T_58458}; // @[Mux.scala 19:72:@32180.4]
  assign _T_58597 = _T_2704 ? _T_58595 : 16'h0; // @[Mux.scala 19:72:@32181.4]
  assign _T_58598 = _T_58342 | _T_58359; // @[Mux.scala 19:72:@32182.4]
  assign _T_58599 = _T_58598 | _T_58376; // @[Mux.scala 19:72:@32183.4]
  assign _T_58600 = _T_58599 | _T_58393; // @[Mux.scala 19:72:@32184.4]
  assign _T_58601 = _T_58600 | _T_58410; // @[Mux.scala 19:72:@32185.4]
  assign _T_58602 = _T_58601 | _T_58427; // @[Mux.scala 19:72:@32186.4]
  assign _T_58603 = _T_58602 | _T_58444; // @[Mux.scala 19:72:@32187.4]
  assign _T_58604 = _T_58603 | _T_58461; // @[Mux.scala 19:72:@32188.4]
  assign _T_58605 = _T_58604 | _T_58478; // @[Mux.scala 19:72:@32189.4]
  assign _T_58606 = _T_58605 | _T_58495; // @[Mux.scala 19:72:@32190.4]
  assign _T_58607 = _T_58606 | _T_58512; // @[Mux.scala 19:72:@32191.4]
  assign _T_58608 = _T_58607 | _T_58529; // @[Mux.scala 19:72:@32192.4]
  assign _T_58609 = _T_58608 | _T_58546; // @[Mux.scala 19:72:@32193.4]
  assign _T_58610 = _T_58609 | _T_58563; // @[Mux.scala 19:72:@32194.4]
  assign _T_58611 = _T_58610 | _T_58580; // @[Mux.scala 19:72:@32195.4]
  assign _T_58612 = _T_58611 | _T_58597; // @[Mux.scala 19:72:@32196.4]
  assign _T_59190 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0}; // @[Mux.scala 19:72:@32546.4]
  assign _T_59197 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8}; // @[Mux.scala 19:72:@32553.4]
  assign _T_59198 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,_T_59190}; // @[Mux.scala 19:72:@32554.4]
  assign _T_59200 = _T_2689 ? _T_59198 : 16'h0; // @[Mux.scala 19:72:@32555.4]
  assign _T_59207 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1}; // @[Mux.scala 19:72:@32562.4]
  assign _T_59214 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9}; // @[Mux.scala 19:72:@32569.4]
  assign _T_59215 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,_T_59207}; // @[Mux.scala 19:72:@32570.4]
  assign _T_59217 = _T_2690 ? _T_59215 : 16'h0; // @[Mux.scala 19:72:@32571.4]
  assign _T_59224 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2}; // @[Mux.scala 19:72:@32578.4]
  assign _T_59231 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10}; // @[Mux.scala 19:72:@32585.4]
  assign _T_59232 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,_T_59224}; // @[Mux.scala 19:72:@32586.4]
  assign _T_59234 = _T_2691 ? _T_59232 : 16'h0; // @[Mux.scala 19:72:@32587.4]
  assign _T_59241 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3}; // @[Mux.scala 19:72:@32594.4]
  assign _T_59248 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11}; // @[Mux.scala 19:72:@32601.4]
  assign _T_59249 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,_T_59241}; // @[Mux.scala 19:72:@32602.4]
  assign _T_59251 = _T_2692 ? _T_59249 : 16'h0; // @[Mux.scala 19:72:@32603.4]
  assign _T_59258 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4}; // @[Mux.scala 19:72:@32610.4]
  assign _T_59265 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12}; // @[Mux.scala 19:72:@32617.4]
  assign _T_59266 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,_T_59258}; // @[Mux.scala 19:72:@32618.4]
  assign _T_59268 = _T_2693 ? _T_59266 : 16'h0; // @[Mux.scala 19:72:@32619.4]
  assign _T_59275 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5}; // @[Mux.scala 19:72:@32626.4]
  assign _T_59282 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13}; // @[Mux.scala 19:72:@32633.4]
  assign _T_59283 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,_T_59275}; // @[Mux.scala 19:72:@32634.4]
  assign _T_59285 = _T_2694 ? _T_59283 : 16'h0; // @[Mux.scala 19:72:@32635.4]
  assign _T_59292 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6}; // @[Mux.scala 19:72:@32642.4]
  assign _T_59299 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14}; // @[Mux.scala 19:72:@32649.4]
  assign _T_59300 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,_T_59292}; // @[Mux.scala 19:72:@32650.4]
  assign _T_59302 = _T_2695 ? _T_59300 : 16'h0; // @[Mux.scala 19:72:@32651.4]
  assign _T_59309 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7}; // @[Mux.scala 19:72:@32658.4]
  assign _T_59316 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15}; // @[Mux.scala 19:72:@32665.4]
  assign _T_59317 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,_T_59309}; // @[Mux.scala 19:72:@32666.4]
  assign _T_59319 = _T_2696 ? _T_59317 : 16'h0; // @[Mux.scala 19:72:@32667.4]
  assign _T_59334 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,_T_59197}; // @[Mux.scala 19:72:@32682.4]
  assign _T_59336 = _T_2697 ? _T_59334 : 16'h0; // @[Mux.scala 19:72:@32683.4]
  assign _T_59351 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,_T_59214}; // @[Mux.scala 19:72:@32698.4]
  assign _T_59353 = _T_2698 ? _T_59351 : 16'h0; // @[Mux.scala 19:72:@32699.4]
  assign _T_59368 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,_T_59231}; // @[Mux.scala 19:72:@32714.4]
  assign _T_59370 = _T_2699 ? _T_59368 : 16'h0; // @[Mux.scala 19:72:@32715.4]
  assign _T_59385 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,_T_59248}; // @[Mux.scala 19:72:@32730.4]
  assign _T_59387 = _T_2700 ? _T_59385 : 16'h0; // @[Mux.scala 19:72:@32731.4]
  assign _T_59402 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,_T_59265}; // @[Mux.scala 19:72:@32746.4]
  assign _T_59404 = _T_2701 ? _T_59402 : 16'h0; // @[Mux.scala 19:72:@32747.4]
  assign _T_59419 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,_T_59282}; // @[Mux.scala 19:72:@32762.4]
  assign _T_59421 = _T_2702 ? _T_59419 : 16'h0; // @[Mux.scala 19:72:@32763.4]
  assign _T_59436 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,_T_59299}; // @[Mux.scala 19:72:@32778.4]
  assign _T_59438 = _T_2703 ? _T_59436 : 16'h0; // @[Mux.scala 19:72:@32779.4]
  assign _T_59453 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,_T_59316}; // @[Mux.scala 19:72:@32794.4]
  assign _T_59455 = _T_2704 ? _T_59453 : 16'h0; // @[Mux.scala 19:72:@32795.4]
  assign _T_59456 = _T_59200 | _T_59217; // @[Mux.scala 19:72:@32796.4]
  assign _T_59457 = _T_59456 | _T_59234; // @[Mux.scala 19:72:@32797.4]
  assign _T_59458 = _T_59457 | _T_59251; // @[Mux.scala 19:72:@32798.4]
  assign _T_59459 = _T_59458 | _T_59268; // @[Mux.scala 19:72:@32799.4]
  assign _T_59460 = _T_59459 | _T_59285; // @[Mux.scala 19:72:@32800.4]
  assign _T_59461 = _T_59460 | _T_59302; // @[Mux.scala 19:72:@32801.4]
  assign _T_59462 = _T_59461 | _T_59319; // @[Mux.scala 19:72:@32802.4]
  assign _T_59463 = _T_59462 | _T_59336; // @[Mux.scala 19:72:@32803.4]
  assign _T_59464 = _T_59463 | _T_59353; // @[Mux.scala 19:72:@32804.4]
  assign _T_59465 = _T_59464 | _T_59370; // @[Mux.scala 19:72:@32805.4]
  assign _T_59466 = _T_59465 | _T_59387; // @[Mux.scala 19:72:@32806.4]
  assign _T_59467 = _T_59466 | _T_59404; // @[Mux.scala 19:72:@32807.4]
  assign _T_59468 = _T_59467 | _T_59421; // @[Mux.scala 19:72:@32808.4]
  assign _T_59469 = _T_59468 | _T_59438; // @[Mux.scala 19:72:@32809.4]
  assign _T_59470 = _T_59469 | _T_59455; // @[Mux.scala 19:72:@32810.4]
  assign _T_60048 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0}; // @[Mux.scala 19:72:@33160.4]
  assign _T_60055 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8}; // @[Mux.scala 19:72:@33167.4]
  assign _T_60056 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,_T_60048}; // @[Mux.scala 19:72:@33168.4]
  assign _T_60058 = _T_2689 ? _T_60056 : 16'h0; // @[Mux.scala 19:72:@33169.4]
  assign _T_60065 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1}; // @[Mux.scala 19:72:@33176.4]
  assign _T_60072 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9}; // @[Mux.scala 19:72:@33183.4]
  assign _T_60073 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,_T_60065}; // @[Mux.scala 19:72:@33184.4]
  assign _T_60075 = _T_2690 ? _T_60073 : 16'h0; // @[Mux.scala 19:72:@33185.4]
  assign _T_60082 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2}; // @[Mux.scala 19:72:@33192.4]
  assign _T_60089 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10}; // @[Mux.scala 19:72:@33199.4]
  assign _T_60090 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,_T_60082}; // @[Mux.scala 19:72:@33200.4]
  assign _T_60092 = _T_2691 ? _T_60090 : 16'h0; // @[Mux.scala 19:72:@33201.4]
  assign _T_60099 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3}; // @[Mux.scala 19:72:@33208.4]
  assign _T_60106 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11}; // @[Mux.scala 19:72:@33215.4]
  assign _T_60107 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,_T_60099}; // @[Mux.scala 19:72:@33216.4]
  assign _T_60109 = _T_2692 ? _T_60107 : 16'h0; // @[Mux.scala 19:72:@33217.4]
  assign _T_60116 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4}; // @[Mux.scala 19:72:@33224.4]
  assign _T_60123 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12}; // @[Mux.scala 19:72:@33231.4]
  assign _T_60124 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,_T_60116}; // @[Mux.scala 19:72:@33232.4]
  assign _T_60126 = _T_2693 ? _T_60124 : 16'h0; // @[Mux.scala 19:72:@33233.4]
  assign _T_60133 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5}; // @[Mux.scala 19:72:@33240.4]
  assign _T_60140 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13}; // @[Mux.scala 19:72:@33247.4]
  assign _T_60141 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,_T_60133}; // @[Mux.scala 19:72:@33248.4]
  assign _T_60143 = _T_2694 ? _T_60141 : 16'h0; // @[Mux.scala 19:72:@33249.4]
  assign _T_60150 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6}; // @[Mux.scala 19:72:@33256.4]
  assign _T_60157 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14}; // @[Mux.scala 19:72:@33263.4]
  assign _T_60158 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,_T_60150}; // @[Mux.scala 19:72:@33264.4]
  assign _T_60160 = _T_2695 ? _T_60158 : 16'h0; // @[Mux.scala 19:72:@33265.4]
  assign _T_60167 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7}; // @[Mux.scala 19:72:@33272.4]
  assign _T_60174 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15}; // @[Mux.scala 19:72:@33279.4]
  assign _T_60175 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,_T_60167}; // @[Mux.scala 19:72:@33280.4]
  assign _T_60177 = _T_2696 ? _T_60175 : 16'h0; // @[Mux.scala 19:72:@33281.4]
  assign _T_60192 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,_T_60055}; // @[Mux.scala 19:72:@33296.4]
  assign _T_60194 = _T_2697 ? _T_60192 : 16'h0; // @[Mux.scala 19:72:@33297.4]
  assign _T_60209 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,_T_60072}; // @[Mux.scala 19:72:@33312.4]
  assign _T_60211 = _T_2698 ? _T_60209 : 16'h0; // @[Mux.scala 19:72:@33313.4]
  assign _T_60226 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,_T_60089}; // @[Mux.scala 19:72:@33328.4]
  assign _T_60228 = _T_2699 ? _T_60226 : 16'h0; // @[Mux.scala 19:72:@33329.4]
  assign _T_60243 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,_T_60106}; // @[Mux.scala 19:72:@33344.4]
  assign _T_60245 = _T_2700 ? _T_60243 : 16'h0; // @[Mux.scala 19:72:@33345.4]
  assign _T_60260 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,_T_60123}; // @[Mux.scala 19:72:@33360.4]
  assign _T_60262 = _T_2701 ? _T_60260 : 16'h0; // @[Mux.scala 19:72:@33361.4]
  assign _T_60277 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,_T_60140}; // @[Mux.scala 19:72:@33376.4]
  assign _T_60279 = _T_2702 ? _T_60277 : 16'h0; // @[Mux.scala 19:72:@33377.4]
  assign _T_60294 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,_T_60157}; // @[Mux.scala 19:72:@33392.4]
  assign _T_60296 = _T_2703 ? _T_60294 : 16'h0; // @[Mux.scala 19:72:@33393.4]
  assign _T_60311 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,_T_60174}; // @[Mux.scala 19:72:@33408.4]
  assign _T_60313 = _T_2704 ? _T_60311 : 16'h0; // @[Mux.scala 19:72:@33409.4]
  assign _T_60314 = _T_60058 | _T_60075; // @[Mux.scala 19:72:@33410.4]
  assign _T_60315 = _T_60314 | _T_60092; // @[Mux.scala 19:72:@33411.4]
  assign _T_60316 = _T_60315 | _T_60109; // @[Mux.scala 19:72:@33412.4]
  assign _T_60317 = _T_60316 | _T_60126; // @[Mux.scala 19:72:@33413.4]
  assign _T_60318 = _T_60317 | _T_60143; // @[Mux.scala 19:72:@33414.4]
  assign _T_60319 = _T_60318 | _T_60160; // @[Mux.scala 19:72:@33415.4]
  assign _T_60320 = _T_60319 | _T_60177; // @[Mux.scala 19:72:@33416.4]
  assign _T_60321 = _T_60320 | _T_60194; // @[Mux.scala 19:72:@33417.4]
  assign _T_60322 = _T_60321 | _T_60211; // @[Mux.scala 19:72:@33418.4]
  assign _T_60323 = _T_60322 | _T_60228; // @[Mux.scala 19:72:@33419.4]
  assign _T_60324 = _T_60323 | _T_60245; // @[Mux.scala 19:72:@33420.4]
  assign _T_60325 = _T_60324 | _T_60262; // @[Mux.scala 19:72:@33421.4]
  assign _T_60326 = _T_60325 | _T_60279; // @[Mux.scala 19:72:@33422.4]
  assign _T_60327 = _T_60326 | _T_60296; // @[Mux.scala 19:72:@33423.4]
  assign _T_60328 = _T_60327 | _T_60313; // @[Mux.scala 19:72:@33424.4]
  assign _T_60906 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0}; // @[Mux.scala 19:72:@33774.4]
  assign _T_60913 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8}; // @[Mux.scala 19:72:@33781.4]
  assign _T_60914 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,_T_60906}; // @[Mux.scala 19:72:@33782.4]
  assign _T_60916 = _T_2689 ? _T_60914 : 16'h0; // @[Mux.scala 19:72:@33783.4]
  assign _T_60923 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1}; // @[Mux.scala 19:72:@33790.4]
  assign _T_60930 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9}; // @[Mux.scala 19:72:@33797.4]
  assign _T_60931 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,_T_60923}; // @[Mux.scala 19:72:@33798.4]
  assign _T_60933 = _T_2690 ? _T_60931 : 16'h0; // @[Mux.scala 19:72:@33799.4]
  assign _T_60940 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2}; // @[Mux.scala 19:72:@33806.4]
  assign _T_60947 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10}; // @[Mux.scala 19:72:@33813.4]
  assign _T_60948 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,_T_60940}; // @[Mux.scala 19:72:@33814.4]
  assign _T_60950 = _T_2691 ? _T_60948 : 16'h0; // @[Mux.scala 19:72:@33815.4]
  assign _T_60957 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3}; // @[Mux.scala 19:72:@33822.4]
  assign _T_60964 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11}; // @[Mux.scala 19:72:@33829.4]
  assign _T_60965 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,_T_60957}; // @[Mux.scala 19:72:@33830.4]
  assign _T_60967 = _T_2692 ? _T_60965 : 16'h0; // @[Mux.scala 19:72:@33831.4]
  assign _T_60974 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4}; // @[Mux.scala 19:72:@33838.4]
  assign _T_60981 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12}; // @[Mux.scala 19:72:@33845.4]
  assign _T_60982 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,_T_60974}; // @[Mux.scala 19:72:@33846.4]
  assign _T_60984 = _T_2693 ? _T_60982 : 16'h0; // @[Mux.scala 19:72:@33847.4]
  assign _T_60991 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5}; // @[Mux.scala 19:72:@33854.4]
  assign _T_60998 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13}; // @[Mux.scala 19:72:@33861.4]
  assign _T_60999 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,_T_60991}; // @[Mux.scala 19:72:@33862.4]
  assign _T_61001 = _T_2694 ? _T_60999 : 16'h0; // @[Mux.scala 19:72:@33863.4]
  assign _T_61008 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6}; // @[Mux.scala 19:72:@33870.4]
  assign _T_61015 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14}; // @[Mux.scala 19:72:@33877.4]
  assign _T_61016 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,_T_61008}; // @[Mux.scala 19:72:@33878.4]
  assign _T_61018 = _T_2695 ? _T_61016 : 16'h0; // @[Mux.scala 19:72:@33879.4]
  assign _T_61025 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7}; // @[Mux.scala 19:72:@33886.4]
  assign _T_61032 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15}; // @[Mux.scala 19:72:@33893.4]
  assign _T_61033 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,_T_61025}; // @[Mux.scala 19:72:@33894.4]
  assign _T_61035 = _T_2696 ? _T_61033 : 16'h0; // @[Mux.scala 19:72:@33895.4]
  assign _T_61050 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,_T_60913}; // @[Mux.scala 19:72:@33910.4]
  assign _T_61052 = _T_2697 ? _T_61050 : 16'h0; // @[Mux.scala 19:72:@33911.4]
  assign _T_61067 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,_T_60930}; // @[Mux.scala 19:72:@33926.4]
  assign _T_61069 = _T_2698 ? _T_61067 : 16'h0; // @[Mux.scala 19:72:@33927.4]
  assign _T_61084 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,_T_60947}; // @[Mux.scala 19:72:@33942.4]
  assign _T_61086 = _T_2699 ? _T_61084 : 16'h0; // @[Mux.scala 19:72:@33943.4]
  assign _T_61101 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,_T_60964}; // @[Mux.scala 19:72:@33958.4]
  assign _T_61103 = _T_2700 ? _T_61101 : 16'h0; // @[Mux.scala 19:72:@33959.4]
  assign _T_61118 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,_T_60981}; // @[Mux.scala 19:72:@33974.4]
  assign _T_61120 = _T_2701 ? _T_61118 : 16'h0; // @[Mux.scala 19:72:@33975.4]
  assign _T_61135 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,_T_60998}; // @[Mux.scala 19:72:@33990.4]
  assign _T_61137 = _T_2702 ? _T_61135 : 16'h0; // @[Mux.scala 19:72:@33991.4]
  assign _T_61152 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,_T_61015}; // @[Mux.scala 19:72:@34006.4]
  assign _T_61154 = _T_2703 ? _T_61152 : 16'h0; // @[Mux.scala 19:72:@34007.4]
  assign _T_61169 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,_T_61032}; // @[Mux.scala 19:72:@34022.4]
  assign _T_61171 = _T_2704 ? _T_61169 : 16'h0; // @[Mux.scala 19:72:@34023.4]
  assign _T_61172 = _T_60916 | _T_60933; // @[Mux.scala 19:72:@34024.4]
  assign _T_61173 = _T_61172 | _T_60950; // @[Mux.scala 19:72:@34025.4]
  assign _T_61174 = _T_61173 | _T_60967; // @[Mux.scala 19:72:@34026.4]
  assign _T_61175 = _T_61174 | _T_60984; // @[Mux.scala 19:72:@34027.4]
  assign _T_61176 = _T_61175 | _T_61001; // @[Mux.scala 19:72:@34028.4]
  assign _T_61177 = _T_61176 | _T_61018; // @[Mux.scala 19:72:@34029.4]
  assign _T_61178 = _T_61177 | _T_61035; // @[Mux.scala 19:72:@34030.4]
  assign _T_61179 = _T_61178 | _T_61052; // @[Mux.scala 19:72:@34031.4]
  assign _T_61180 = _T_61179 | _T_61069; // @[Mux.scala 19:72:@34032.4]
  assign _T_61181 = _T_61180 | _T_61086; // @[Mux.scala 19:72:@34033.4]
  assign _T_61182 = _T_61181 | _T_61103; // @[Mux.scala 19:72:@34034.4]
  assign _T_61183 = _T_61182 | _T_61120; // @[Mux.scala 19:72:@34035.4]
  assign _T_61184 = _T_61183 | _T_61137; // @[Mux.scala 19:72:@34036.4]
  assign _T_61185 = _T_61184 | _T_61154; // @[Mux.scala 19:72:@34037.4]
  assign _T_61186 = _T_61185 | _T_61171; // @[Mux.scala 19:72:@34038.4]
  assign _T_61764 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0}; // @[Mux.scala 19:72:@34388.4]
  assign _T_61771 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8}; // @[Mux.scala 19:72:@34395.4]
  assign _T_61772 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,_T_61764}; // @[Mux.scala 19:72:@34396.4]
  assign _T_61774 = _T_2689 ? _T_61772 : 16'h0; // @[Mux.scala 19:72:@34397.4]
  assign _T_61781 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1}; // @[Mux.scala 19:72:@34404.4]
  assign _T_61788 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9}; // @[Mux.scala 19:72:@34411.4]
  assign _T_61789 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,_T_61781}; // @[Mux.scala 19:72:@34412.4]
  assign _T_61791 = _T_2690 ? _T_61789 : 16'h0; // @[Mux.scala 19:72:@34413.4]
  assign _T_61798 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2}; // @[Mux.scala 19:72:@34420.4]
  assign _T_61805 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10}; // @[Mux.scala 19:72:@34427.4]
  assign _T_61806 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,_T_61798}; // @[Mux.scala 19:72:@34428.4]
  assign _T_61808 = _T_2691 ? _T_61806 : 16'h0; // @[Mux.scala 19:72:@34429.4]
  assign _T_61815 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3}; // @[Mux.scala 19:72:@34436.4]
  assign _T_61822 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11}; // @[Mux.scala 19:72:@34443.4]
  assign _T_61823 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,_T_61815}; // @[Mux.scala 19:72:@34444.4]
  assign _T_61825 = _T_2692 ? _T_61823 : 16'h0; // @[Mux.scala 19:72:@34445.4]
  assign _T_61832 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4}; // @[Mux.scala 19:72:@34452.4]
  assign _T_61839 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12}; // @[Mux.scala 19:72:@34459.4]
  assign _T_61840 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,_T_61832}; // @[Mux.scala 19:72:@34460.4]
  assign _T_61842 = _T_2693 ? _T_61840 : 16'h0; // @[Mux.scala 19:72:@34461.4]
  assign _T_61849 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5}; // @[Mux.scala 19:72:@34468.4]
  assign _T_61856 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13}; // @[Mux.scala 19:72:@34475.4]
  assign _T_61857 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,_T_61849}; // @[Mux.scala 19:72:@34476.4]
  assign _T_61859 = _T_2694 ? _T_61857 : 16'h0; // @[Mux.scala 19:72:@34477.4]
  assign _T_61866 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6}; // @[Mux.scala 19:72:@34484.4]
  assign _T_61873 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14}; // @[Mux.scala 19:72:@34491.4]
  assign _T_61874 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,_T_61866}; // @[Mux.scala 19:72:@34492.4]
  assign _T_61876 = _T_2695 ? _T_61874 : 16'h0; // @[Mux.scala 19:72:@34493.4]
  assign _T_61883 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7}; // @[Mux.scala 19:72:@34500.4]
  assign _T_61890 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15}; // @[Mux.scala 19:72:@34507.4]
  assign _T_61891 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,_T_61883}; // @[Mux.scala 19:72:@34508.4]
  assign _T_61893 = _T_2696 ? _T_61891 : 16'h0; // @[Mux.scala 19:72:@34509.4]
  assign _T_61908 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,_T_61771}; // @[Mux.scala 19:72:@34524.4]
  assign _T_61910 = _T_2697 ? _T_61908 : 16'h0; // @[Mux.scala 19:72:@34525.4]
  assign _T_61925 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,_T_61788}; // @[Mux.scala 19:72:@34540.4]
  assign _T_61927 = _T_2698 ? _T_61925 : 16'h0; // @[Mux.scala 19:72:@34541.4]
  assign _T_61942 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,_T_61805}; // @[Mux.scala 19:72:@34556.4]
  assign _T_61944 = _T_2699 ? _T_61942 : 16'h0; // @[Mux.scala 19:72:@34557.4]
  assign _T_61959 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,_T_61822}; // @[Mux.scala 19:72:@34572.4]
  assign _T_61961 = _T_2700 ? _T_61959 : 16'h0; // @[Mux.scala 19:72:@34573.4]
  assign _T_61976 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,_T_61839}; // @[Mux.scala 19:72:@34588.4]
  assign _T_61978 = _T_2701 ? _T_61976 : 16'h0; // @[Mux.scala 19:72:@34589.4]
  assign _T_61993 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,_T_61856}; // @[Mux.scala 19:72:@34604.4]
  assign _T_61995 = _T_2702 ? _T_61993 : 16'h0; // @[Mux.scala 19:72:@34605.4]
  assign _T_62010 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,_T_61873}; // @[Mux.scala 19:72:@34620.4]
  assign _T_62012 = _T_2703 ? _T_62010 : 16'h0; // @[Mux.scala 19:72:@34621.4]
  assign _T_62027 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,_T_61890}; // @[Mux.scala 19:72:@34636.4]
  assign _T_62029 = _T_2704 ? _T_62027 : 16'h0; // @[Mux.scala 19:72:@34637.4]
  assign _T_62030 = _T_61774 | _T_61791; // @[Mux.scala 19:72:@34638.4]
  assign _T_62031 = _T_62030 | _T_61808; // @[Mux.scala 19:72:@34639.4]
  assign _T_62032 = _T_62031 | _T_61825; // @[Mux.scala 19:72:@34640.4]
  assign _T_62033 = _T_62032 | _T_61842; // @[Mux.scala 19:72:@34641.4]
  assign _T_62034 = _T_62033 | _T_61859; // @[Mux.scala 19:72:@34642.4]
  assign _T_62035 = _T_62034 | _T_61876; // @[Mux.scala 19:72:@34643.4]
  assign _T_62036 = _T_62035 | _T_61893; // @[Mux.scala 19:72:@34644.4]
  assign _T_62037 = _T_62036 | _T_61910; // @[Mux.scala 19:72:@34645.4]
  assign _T_62038 = _T_62037 | _T_61927; // @[Mux.scala 19:72:@34646.4]
  assign _T_62039 = _T_62038 | _T_61944; // @[Mux.scala 19:72:@34647.4]
  assign _T_62040 = _T_62039 | _T_61961; // @[Mux.scala 19:72:@34648.4]
  assign _T_62041 = _T_62040 | _T_61978; // @[Mux.scala 19:72:@34649.4]
  assign _T_62042 = _T_62041 | _T_61995; // @[Mux.scala 19:72:@34650.4]
  assign _T_62043 = _T_62042 | _T_62012; // @[Mux.scala 19:72:@34651.4]
  assign _T_62044 = _T_62043 | _T_62029; // @[Mux.scala 19:72:@34652.4]
  assign _T_62622 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0}; // @[Mux.scala 19:72:@35002.4]
  assign _T_62629 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8}; // @[Mux.scala 19:72:@35009.4]
  assign _T_62630 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,_T_62622}; // @[Mux.scala 19:72:@35010.4]
  assign _T_62632 = _T_2689 ? _T_62630 : 16'h0; // @[Mux.scala 19:72:@35011.4]
  assign _T_62639 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1}; // @[Mux.scala 19:72:@35018.4]
  assign _T_62646 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9}; // @[Mux.scala 19:72:@35025.4]
  assign _T_62647 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,_T_62639}; // @[Mux.scala 19:72:@35026.4]
  assign _T_62649 = _T_2690 ? _T_62647 : 16'h0; // @[Mux.scala 19:72:@35027.4]
  assign _T_62656 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2}; // @[Mux.scala 19:72:@35034.4]
  assign _T_62663 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10}; // @[Mux.scala 19:72:@35041.4]
  assign _T_62664 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,_T_62656}; // @[Mux.scala 19:72:@35042.4]
  assign _T_62666 = _T_2691 ? _T_62664 : 16'h0; // @[Mux.scala 19:72:@35043.4]
  assign _T_62673 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3}; // @[Mux.scala 19:72:@35050.4]
  assign _T_62680 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11}; // @[Mux.scala 19:72:@35057.4]
  assign _T_62681 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,_T_62673}; // @[Mux.scala 19:72:@35058.4]
  assign _T_62683 = _T_2692 ? _T_62681 : 16'h0; // @[Mux.scala 19:72:@35059.4]
  assign _T_62690 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4}; // @[Mux.scala 19:72:@35066.4]
  assign _T_62697 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12}; // @[Mux.scala 19:72:@35073.4]
  assign _T_62698 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,_T_62690}; // @[Mux.scala 19:72:@35074.4]
  assign _T_62700 = _T_2693 ? _T_62698 : 16'h0; // @[Mux.scala 19:72:@35075.4]
  assign _T_62707 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5}; // @[Mux.scala 19:72:@35082.4]
  assign _T_62714 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13}; // @[Mux.scala 19:72:@35089.4]
  assign _T_62715 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,_T_62707}; // @[Mux.scala 19:72:@35090.4]
  assign _T_62717 = _T_2694 ? _T_62715 : 16'h0; // @[Mux.scala 19:72:@35091.4]
  assign _T_62724 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6}; // @[Mux.scala 19:72:@35098.4]
  assign _T_62731 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14}; // @[Mux.scala 19:72:@35105.4]
  assign _T_62732 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,_T_62724}; // @[Mux.scala 19:72:@35106.4]
  assign _T_62734 = _T_2695 ? _T_62732 : 16'h0; // @[Mux.scala 19:72:@35107.4]
  assign _T_62741 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7}; // @[Mux.scala 19:72:@35114.4]
  assign _T_62748 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15}; // @[Mux.scala 19:72:@35121.4]
  assign _T_62749 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,_T_62741}; // @[Mux.scala 19:72:@35122.4]
  assign _T_62751 = _T_2696 ? _T_62749 : 16'h0; // @[Mux.scala 19:72:@35123.4]
  assign _T_62766 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,_T_62629}; // @[Mux.scala 19:72:@35138.4]
  assign _T_62768 = _T_2697 ? _T_62766 : 16'h0; // @[Mux.scala 19:72:@35139.4]
  assign _T_62783 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,_T_62646}; // @[Mux.scala 19:72:@35154.4]
  assign _T_62785 = _T_2698 ? _T_62783 : 16'h0; // @[Mux.scala 19:72:@35155.4]
  assign _T_62800 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,_T_62663}; // @[Mux.scala 19:72:@35170.4]
  assign _T_62802 = _T_2699 ? _T_62800 : 16'h0; // @[Mux.scala 19:72:@35171.4]
  assign _T_62817 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,_T_62680}; // @[Mux.scala 19:72:@35186.4]
  assign _T_62819 = _T_2700 ? _T_62817 : 16'h0; // @[Mux.scala 19:72:@35187.4]
  assign _T_62834 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,_T_62697}; // @[Mux.scala 19:72:@35202.4]
  assign _T_62836 = _T_2701 ? _T_62834 : 16'h0; // @[Mux.scala 19:72:@35203.4]
  assign _T_62851 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,_T_62714}; // @[Mux.scala 19:72:@35218.4]
  assign _T_62853 = _T_2702 ? _T_62851 : 16'h0; // @[Mux.scala 19:72:@35219.4]
  assign _T_62868 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,_T_62731}; // @[Mux.scala 19:72:@35234.4]
  assign _T_62870 = _T_2703 ? _T_62868 : 16'h0; // @[Mux.scala 19:72:@35235.4]
  assign _T_62885 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,_T_62748}; // @[Mux.scala 19:72:@35250.4]
  assign _T_62887 = _T_2704 ? _T_62885 : 16'h0; // @[Mux.scala 19:72:@35251.4]
  assign _T_62888 = _T_62632 | _T_62649; // @[Mux.scala 19:72:@35252.4]
  assign _T_62889 = _T_62888 | _T_62666; // @[Mux.scala 19:72:@35253.4]
  assign _T_62890 = _T_62889 | _T_62683; // @[Mux.scala 19:72:@35254.4]
  assign _T_62891 = _T_62890 | _T_62700; // @[Mux.scala 19:72:@35255.4]
  assign _T_62892 = _T_62891 | _T_62717; // @[Mux.scala 19:72:@35256.4]
  assign _T_62893 = _T_62892 | _T_62734; // @[Mux.scala 19:72:@35257.4]
  assign _T_62894 = _T_62893 | _T_62751; // @[Mux.scala 19:72:@35258.4]
  assign _T_62895 = _T_62894 | _T_62768; // @[Mux.scala 19:72:@35259.4]
  assign _T_62896 = _T_62895 | _T_62785; // @[Mux.scala 19:72:@35260.4]
  assign _T_62897 = _T_62896 | _T_62802; // @[Mux.scala 19:72:@35261.4]
  assign _T_62898 = _T_62897 | _T_62819; // @[Mux.scala 19:72:@35262.4]
  assign _T_62899 = _T_62898 | _T_62836; // @[Mux.scala 19:72:@35263.4]
  assign _T_62900 = _T_62899 | _T_62853; // @[Mux.scala 19:72:@35264.4]
  assign _T_62901 = _T_62900 | _T_62870; // @[Mux.scala 19:72:@35265.4]
  assign _T_62902 = _T_62901 | _T_62887; // @[Mux.scala 19:72:@35266.4]
  assign _T_63480 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0}; // @[Mux.scala 19:72:@35616.4]
  assign _T_63487 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8}; // @[Mux.scala 19:72:@35623.4]
  assign _T_63488 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,_T_63480}; // @[Mux.scala 19:72:@35624.4]
  assign _T_63490 = _T_2689 ? _T_63488 : 16'h0; // @[Mux.scala 19:72:@35625.4]
  assign _T_63497 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1}; // @[Mux.scala 19:72:@35632.4]
  assign _T_63504 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9}; // @[Mux.scala 19:72:@35639.4]
  assign _T_63505 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,_T_63497}; // @[Mux.scala 19:72:@35640.4]
  assign _T_63507 = _T_2690 ? _T_63505 : 16'h0; // @[Mux.scala 19:72:@35641.4]
  assign _T_63514 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2}; // @[Mux.scala 19:72:@35648.4]
  assign _T_63521 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10}; // @[Mux.scala 19:72:@35655.4]
  assign _T_63522 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,_T_63514}; // @[Mux.scala 19:72:@35656.4]
  assign _T_63524 = _T_2691 ? _T_63522 : 16'h0; // @[Mux.scala 19:72:@35657.4]
  assign _T_63531 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3}; // @[Mux.scala 19:72:@35664.4]
  assign _T_63538 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11}; // @[Mux.scala 19:72:@35671.4]
  assign _T_63539 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,_T_63531}; // @[Mux.scala 19:72:@35672.4]
  assign _T_63541 = _T_2692 ? _T_63539 : 16'h0; // @[Mux.scala 19:72:@35673.4]
  assign _T_63548 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4}; // @[Mux.scala 19:72:@35680.4]
  assign _T_63555 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12}; // @[Mux.scala 19:72:@35687.4]
  assign _T_63556 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,_T_63548}; // @[Mux.scala 19:72:@35688.4]
  assign _T_63558 = _T_2693 ? _T_63556 : 16'h0; // @[Mux.scala 19:72:@35689.4]
  assign _T_63565 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5}; // @[Mux.scala 19:72:@35696.4]
  assign _T_63572 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13}; // @[Mux.scala 19:72:@35703.4]
  assign _T_63573 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,_T_63565}; // @[Mux.scala 19:72:@35704.4]
  assign _T_63575 = _T_2694 ? _T_63573 : 16'h0; // @[Mux.scala 19:72:@35705.4]
  assign _T_63582 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6}; // @[Mux.scala 19:72:@35712.4]
  assign _T_63589 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14}; // @[Mux.scala 19:72:@35719.4]
  assign _T_63590 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,_T_63582}; // @[Mux.scala 19:72:@35720.4]
  assign _T_63592 = _T_2695 ? _T_63590 : 16'h0; // @[Mux.scala 19:72:@35721.4]
  assign _T_63599 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7}; // @[Mux.scala 19:72:@35728.4]
  assign _T_63606 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15}; // @[Mux.scala 19:72:@35735.4]
  assign _T_63607 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,_T_63599}; // @[Mux.scala 19:72:@35736.4]
  assign _T_63609 = _T_2696 ? _T_63607 : 16'h0; // @[Mux.scala 19:72:@35737.4]
  assign _T_63624 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,_T_63487}; // @[Mux.scala 19:72:@35752.4]
  assign _T_63626 = _T_2697 ? _T_63624 : 16'h0; // @[Mux.scala 19:72:@35753.4]
  assign _T_63641 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,_T_63504}; // @[Mux.scala 19:72:@35768.4]
  assign _T_63643 = _T_2698 ? _T_63641 : 16'h0; // @[Mux.scala 19:72:@35769.4]
  assign _T_63658 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,_T_63521}; // @[Mux.scala 19:72:@35784.4]
  assign _T_63660 = _T_2699 ? _T_63658 : 16'h0; // @[Mux.scala 19:72:@35785.4]
  assign _T_63675 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,_T_63538}; // @[Mux.scala 19:72:@35800.4]
  assign _T_63677 = _T_2700 ? _T_63675 : 16'h0; // @[Mux.scala 19:72:@35801.4]
  assign _T_63692 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,_T_63555}; // @[Mux.scala 19:72:@35816.4]
  assign _T_63694 = _T_2701 ? _T_63692 : 16'h0; // @[Mux.scala 19:72:@35817.4]
  assign _T_63709 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,_T_63572}; // @[Mux.scala 19:72:@35832.4]
  assign _T_63711 = _T_2702 ? _T_63709 : 16'h0; // @[Mux.scala 19:72:@35833.4]
  assign _T_63726 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,_T_63589}; // @[Mux.scala 19:72:@35848.4]
  assign _T_63728 = _T_2703 ? _T_63726 : 16'h0; // @[Mux.scala 19:72:@35849.4]
  assign _T_63743 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,_T_63606}; // @[Mux.scala 19:72:@35864.4]
  assign _T_63745 = _T_2704 ? _T_63743 : 16'h0; // @[Mux.scala 19:72:@35865.4]
  assign _T_63746 = _T_63490 | _T_63507; // @[Mux.scala 19:72:@35866.4]
  assign _T_63747 = _T_63746 | _T_63524; // @[Mux.scala 19:72:@35867.4]
  assign _T_63748 = _T_63747 | _T_63541; // @[Mux.scala 19:72:@35868.4]
  assign _T_63749 = _T_63748 | _T_63558; // @[Mux.scala 19:72:@35869.4]
  assign _T_63750 = _T_63749 | _T_63575; // @[Mux.scala 19:72:@35870.4]
  assign _T_63751 = _T_63750 | _T_63592; // @[Mux.scala 19:72:@35871.4]
  assign _T_63752 = _T_63751 | _T_63609; // @[Mux.scala 19:72:@35872.4]
  assign _T_63753 = _T_63752 | _T_63626; // @[Mux.scala 19:72:@35873.4]
  assign _T_63754 = _T_63753 | _T_63643; // @[Mux.scala 19:72:@35874.4]
  assign _T_63755 = _T_63754 | _T_63660; // @[Mux.scala 19:72:@35875.4]
  assign _T_63756 = _T_63755 | _T_63677; // @[Mux.scala 19:72:@35876.4]
  assign _T_63757 = _T_63756 | _T_63694; // @[Mux.scala 19:72:@35877.4]
  assign _T_63758 = _T_63757 | _T_63711; // @[Mux.scala 19:72:@35878.4]
  assign _T_63759 = _T_63758 | _T_63728; // @[Mux.scala 19:72:@35879.4]
  assign _T_63760 = _T_63759 | _T_63745; // @[Mux.scala 19:72:@35880.4]
  assign _T_64338 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0}; // @[Mux.scala 19:72:@36230.4]
  assign _T_64345 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8}; // @[Mux.scala 19:72:@36237.4]
  assign _T_64346 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,_T_64338}; // @[Mux.scala 19:72:@36238.4]
  assign _T_64348 = _T_2689 ? _T_64346 : 16'h0; // @[Mux.scala 19:72:@36239.4]
  assign _T_64355 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1}; // @[Mux.scala 19:72:@36246.4]
  assign _T_64362 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9}; // @[Mux.scala 19:72:@36253.4]
  assign _T_64363 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,_T_64355}; // @[Mux.scala 19:72:@36254.4]
  assign _T_64365 = _T_2690 ? _T_64363 : 16'h0; // @[Mux.scala 19:72:@36255.4]
  assign _T_64372 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2}; // @[Mux.scala 19:72:@36262.4]
  assign _T_64379 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10}; // @[Mux.scala 19:72:@36269.4]
  assign _T_64380 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,_T_64372}; // @[Mux.scala 19:72:@36270.4]
  assign _T_64382 = _T_2691 ? _T_64380 : 16'h0; // @[Mux.scala 19:72:@36271.4]
  assign _T_64389 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3}; // @[Mux.scala 19:72:@36278.4]
  assign _T_64396 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11}; // @[Mux.scala 19:72:@36285.4]
  assign _T_64397 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,_T_64389}; // @[Mux.scala 19:72:@36286.4]
  assign _T_64399 = _T_2692 ? _T_64397 : 16'h0; // @[Mux.scala 19:72:@36287.4]
  assign _T_64406 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4}; // @[Mux.scala 19:72:@36294.4]
  assign _T_64413 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12}; // @[Mux.scala 19:72:@36301.4]
  assign _T_64414 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,_T_64406}; // @[Mux.scala 19:72:@36302.4]
  assign _T_64416 = _T_2693 ? _T_64414 : 16'h0; // @[Mux.scala 19:72:@36303.4]
  assign _T_64423 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5}; // @[Mux.scala 19:72:@36310.4]
  assign _T_64430 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13}; // @[Mux.scala 19:72:@36317.4]
  assign _T_64431 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,_T_64423}; // @[Mux.scala 19:72:@36318.4]
  assign _T_64433 = _T_2694 ? _T_64431 : 16'h0; // @[Mux.scala 19:72:@36319.4]
  assign _T_64440 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6}; // @[Mux.scala 19:72:@36326.4]
  assign _T_64447 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14}; // @[Mux.scala 19:72:@36333.4]
  assign _T_64448 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,_T_64440}; // @[Mux.scala 19:72:@36334.4]
  assign _T_64450 = _T_2695 ? _T_64448 : 16'h0; // @[Mux.scala 19:72:@36335.4]
  assign _T_64457 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7}; // @[Mux.scala 19:72:@36342.4]
  assign _T_64464 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15}; // @[Mux.scala 19:72:@36349.4]
  assign _T_64465 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,_T_64457}; // @[Mux.scala 19:72:@36350.4]
  assign _T_64467 = _T_2696 ? _T_64465 : 16'h0; // @[Mux.scala 19:72:@36351.4]
  assign _T_64482 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,_T_64345}; // @[Mux.scala 19:72:@36366.4]
  assign _T_64484 = _T_2697 ? _T_64482 : 16'h0; // @[Mux.scala 19:72:@36367.4]
  assign _T_64499 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,_T_64362}; // @[Mux.scala 19:72:@36382.4]
  assign _T_64501 = _T_2698 ? _T_64499 : 16'h0; // @[Mux.scala 19:72:@36383.4]
  assign _T_64516 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,_T_64379}; // @[Mux.scala 19:72:@36398.4]
  assign _T_64518 = _T_2699 ? _T_64516 : 16'h0; // @[Mux.scala 19:72:@36399.4]
  assign _T_64533 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,_T_64396}; // @[Mux.scala 19:72:@36414.4]
  assign _T_64535 = _T_2700 ? _T_64533 : 16'h0; // @[Mux.scala 19:72:@36415.4]
  assign _T_64550 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,_T_64413}; // @[Mux.scala 19:72:@36430.4]
  assign _T_64552 = _T_2701 ? _T_64550 : 16'h0; // @[Mux.scala 19:72:@36431.4]
  assign _T_64567 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,_T_64430}; // @[Mux.scala 19:72:@36446.4]
  assign _T_64569 = _T_2702 ? _T_64567 : 16'h0; // @[Mux.scala 19:72:@36447.4]
  assign _T_64584 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,_T_64447}; // @[Mux.scala 19:72:@36462.4]
  assign _T_64586 = _T_2703 ? _T_64584 : 16'h0; // @[Mux.scala 19:72:@36463.4]
  assign _T_64601 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,_T_64464}; // @[Mux.scala 19:72:@36478.4]
  assign _T_64603 = _T_2704 ? _T_64601 : 16'h0; // @[Mux.scala 19:72:@36479.4]
  assign _T_64604 = _T_64348 | _T_64365; // @[Mux.scala 19:72:@36480.4]
  assign _T_64605 = _T_64604 | _T_64382; // @[Mux.scala 19:72:@36481.4]
  assign _T_64606 = _T_64605 | _T_64399; // @[Mux.scala 19:72:@36482.4]
  assign _T_64607 = _T_64606 | _T_64416; // @[Mux.scala 19:72:@36483.4]
  assign _T_64608 = _T_64607 | _T_64433; // @[Mux.scala 19:72:@36484.4]
  assign _T_64609 = _T_64608 | _T_64450; // @[Mux.scala 19:72:@36485.4]
  assign _T_64610 = _T_64609 | _T_64467; // @[Mux.scala 19:72:@36486.4]
  assign _T_64611 = _T_64610 | _T_64484; // @[Mux.scala 19:72:@36487.4]
  assign _T_64612 = _T_64611 | _T_64501; // @[Mux.scala 19:72:@36488.4]
  assign _T_64613 = _T_64612 | _T_64518; // @[Mux.scala 19:72:@36489.4]
  assign _T_64614 = _T_64613 | _T_64535; // @[Mux.scala 19:72:@36490.4]
  assign _T_64615 = _T_64614 | _T_64552; // @[Mux.scala 19:72:@36491.4]
  assign _T_64616 = _T_64615 | _T_64569; // @[Mux.scala 19:72:@36492.4]
  assign _T_64617 = _T_64616 | _T_64586; // @[Mux.scala 19:72:@36493.4]
  assign _T_64618 = _T_64617 | _T_64603; // @[Mux.scala 19:72:@36494.4]
  assign _T_65196 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0}; // @[Mux.scala 19:72:@36844.4]
  assign _T_65203 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8}; // @[Mux.scala 19:72:@36851.4]
  assign _T_65204 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,_T_65196}; // @[Mux.scala 19:72:@36852.4]
  assign _T_65206 = _T_2689 ? _T_65204 : 16'h0; // @[Mux.scala 19:72:@36853.4]
  assign _T_65213 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1}; // @[Mux.scala 19:72:@36860.4]
  assign _T_65220 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9}; // @[Mux.scala 19:72:@36867.4]
  assign _T_65221 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,_T_65213}; // @[Mux.scala 19:72:@36868.4]
  assign _T_65223 = _T_2690 ? _T_65221 : 16'h0; // @[Mux.scala 19:72:@36869.4]
  assign _T_65230 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2}; // @[Mux.scala 19:72:@36876.4]
  assign _T_65237 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10}; // @[Mux.scala 19:72:@36883.4]
  assign _T_65238 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,_T_65230}; // @[Mux.scala 19:72:@36884.4]
  assign _T_65240 = _T_2691 ? _T_65238 : 16'h0; // @[Mux.scala 19:72:@36885.4]
  assign _T_65247 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3}; // @[Mux.scala 19:72:@36892.4]
  assign _T_65254 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11}; // @[Mux.scala 19:72:@36899.4]
  assign _T_65255 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,_T_65247}; // @[Mux.scala 19:72:@36900.4]
  assign _T_65257 = _T_2692 ? _T_65255 : 16'h0; // @[Mux.scala 19:72:@36901.4]
  assign _T_65264 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4}; // @[Mux.scala 19:72:@36908.4]
  assign _T_65271 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12}; // @[Mux.scala 19:72:@36915.4]
  assign _T_65272 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,_T_65264}; // @[Mux.scala 19:72:@36916.4]
  assign _T_65274 = _T_2693 ? _T_65272 : 16'h0; // @[Mux.scala 19:72:@36917.4]
  assign _T_65281 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5}; // @[Mux.scala 19:72:@36924.4]
  assign _T_65288 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13}; // @[Mux.scala 19:72:@36931.4]
  assign _T_65289 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,_T_65281}; // @[Mux.scala 19:72:@36932.4]
  assign _T_65291 = _T_2694 ? _T_65289 : 16'h0; // @[Mux.scala 19:72:@36933.4]
  assign _T_65298 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6}; // @[Mux.scala 19:72:@36940.4]
  assign _T_65305 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14}; // @[Mux.scala 19:72:@36947.4]
  assign _T_65306 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,_T_65298}; // @[Mux.scala 19:72:@36948.4]
  assign _T_65308 = _T_2695 ? _T_65306 : 16'h0; // @[Mux.scala 19:72:@36949.4]
  assign _T_65315 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7}; // @[Mux.scala 19:72:@36956.4]
  assign _T_65322 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15}; // @[Mux.scala 19:72:@36963.4]
  assign _T_65323 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,_T_65315}; // @[Mux.scala 19:72:@36964.4]
  assign _T_65325 = _T_2696 ? _T_65323 : 16'h0; // @[Mux.scala 19:72:@36965.4]
  assign _T_65340 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,_T_65203}; // @[Mux.scala 19:72:@36980.4]
  assign _T_65342 = _T_2697 ? _T_65340 : 16'h0; // @[Mux.scala 19:72:@36981.4]
  assign _T_65357 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,_T_65220}; // @[Mux.scala 19:72:@36996.4]
  assign _T_65359 = _T_2698 ? _T_65357 : 16'h0; // @[Mux.scala 19:72:@36997.4]
  assign _T_65374 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,_T_65237}; // @[Mux.scala 19:72:@37012.4]
  assign _T_65376 = _T_2699 ? _T_65374 : 16'h0; // @[Mux.scala 19:72:@37013.4]
  assign _T_65391 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,_T_65254}; // @[Mux.scala 19:72:@37028.4]
  assign _T_65393 = _T_2700 ? _T_65391 : 16'h0; // @[Mux.scala 19:72:@37029.4]
  assign _T_65408 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,_T_65271}; // @[Mux.scala 19:72:@37044.4]
  assign _T_65410 = _T_2701 ? _T_65408 : 16'h0; // @[Mux.scala 19:72:@37045.4]
  assign _T_65425 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,_T_65288}; // @[Mux.scala 19:72:@37060.4]
  assign _T_65427 = _T_2702 ? _T_65425 : 16'h0; // @[Mux.scala 19:72:@37061.4]
  assign _T_65442 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,_T_65305}; // @[Mux.scala 19:72:@37076.4]
  assign _T_65444 = _T_2703 ? _T_65442 : 16'h0; // @[Mux.scala 19:72:@37077.4]
  assign _T_65459 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,_T_65322}; // @[Mux.scala 19:72:@37092.4]
  assign _T_65461 = _T_2704 ? _T_65459 : 16'h0; // @[Mux.scala 19:72:@37093.4]
  assign _T_65462 = _T_65206 | _T_65223; // @[Mux.scala 19:72:@37094.4]
  assign _T_65463 = _T_65462 | _T_65240; // @[Mux.scala 19:72:@37095.4]
  assign _T_65464 = _T_65463 | _T_65257; // @[Mux.scala 19:72:@37096.4]
  assign _T_65465 = _T_65464 | _T_65274; // @[Mux.scala 19:72:@37097.4]
  assign _T_65466 = _T_65465 | _T_65291; // @[Mux.scala 19:72:@37098.4]
  assign _T_65467 = _T_65466 | _T_65308; // @[Mux.scala 19:72:@37099.4]
  assign _T_65468 = _T_65467 | _T_65325; // @[Mux.scala 19:72:@37100.4]
  assign _T_65469 = _T_65468 | _T_65342; // @[Mux.scala 19:72:@37101.4]
  assign _T_65470 = _T_65469 | _T_65359; // @[Mux.scala 19:72:@37102.4]
  assign _T_65471 = _T_65470 | _T_65376; // @[Mux.scala 19:72:@37103.4]
  assign _T_65472 = _T_65471 | _T_65393; // @[Mux.scala 19:72:@37104.4]
  assign _T_65473 = _T_65472 | _T_65410; // @[Mux.scala 19:72:@37105.4]
  assign _T_65474 = _T_65473 | _T_65427; // @[Mux.scala 19:72:@37106.4]
  assign _T_65475 = _T_65474 | _T_65444; // @[Mux.scala 19:72:@37107.4]
  assign _T_65476 = _T_65475 | _T_65461; // @[Mux.scala 19:72:@37108.4]
  assign _T_88268 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[LoadQueue.scala 191:60:@37781.4]
  assign _T_88269 = conflictPReg_0_3 ? 2'h3 : _T_88268; // @[LoadQueue.scala 191:60:@37782.4]
  assign _T_88270 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_88269}; // @[LoadQueue.scala 191:60:@37783.4]
  assign _T_88271 = conflictPReg_0_5 ? 3'h5 : _T_88270; // @[LoadQueue.scala 191:60:@37784.4]
  assign _T_88272 = conflictPReg_0_6 ? 3'h6 : _T_88271; // @[LoadQueue.scala 191:60:@37785.4]
  assign _T_88273 = conflictPReg_0_7 ? 3'h7 : _T_88272; // @[LoadQueue.scala 191:60:@37786.4]
  assign _T_88274 = conflictPReg_0_8 ? 4'h8 : {{1'd0}, _T_88273}; // @[LoadQueue.scala 191:60:@37787.4]
  assign _T_88275 = conflictPReg_0_9 ? 4'h9 : _T_88274; // @[LoadQueue.scala 191:60:@37788.4]
  assign _T_88276 = conflictPReg_0_10 ? 4'ha : _T_88275; // @[LoadQueue.scala 191:60:@37789.4]
  assign _T_88277 = conflictPReg_0_11 ? 4'hb : _T_88276; // @[LoadQueue.scala 191:60:@37790.4]
  assign _T_88278 = conflictPReg_0_12 ? 4'hc : _T_88277; // @[LoadQueue.scala 191:60:@37791.4]
  assign _T_88279 = conflictPReg_0_13 ? 4'hd : _T_88278; // @[LoadQueue.scala 191:60:@37792.4]
  assign _T_88280 = conflictPReg_0_14 ? 4'he : _T_88279; // @[LoadQueue.scala 191:60:@37793.4]
  assign _T_88281 = conflictPReg_0_15 ? 4'hf : _T_88280; // @[LoadQueue.scala 191:60:@37794.4]
  assign _T_88284 = conflictPReg_0_0 | conflictPReg_0_1; // @[LoadQueue.scala 192:43:@37796.4]
  assign _T_88285 = _T_88284 | conflictPReg_0_2; // @[LoadQueue.scala 192:43:@37797.4]
  assign _T_88286 = _T_88285 | conflictPReg_0_3; // @[LoadQueue.scala 192:43:@37798.4]
  assign _T_88287 = _T_88286 | conflictPReg_0_4; // @[LoadQueue.scala 192:43:@37799.4]
  assign _T_88288 = _T_88287 | conflictPReg_0_5; // @[LoadQueue.scala 192:43:@37800.4]
  assign _T_88289 = _T_88288 | conflictPReg_0_6; // @[LoadQueue.scala 192:43:@37801.4]
  assign _T_88290 = _T_88289 | conflictPReg_0_7; // @[LoadQueue.scala 192:43:@37802.4]
  assign _T_88291 = _T_88290 | conflictPReg_0_8; // @[LoadQueue.scala 192:43:@37803.4]
  assign _T_88292 = _T_88291 | conflictPReg_0_9; // @[LoadQueue.scala 192:43:@37804.4]
  assign _T_88293 = _T_88292 | conflictPReg_0_10; // @[LoadQueue.scala 192:43:@37805.4]
  assign _T_88294 = _T_88293 | conflictPReg_0_11; // @[LoadQueue.scala 192:43:@37806.4]
  assign _T_88295 = _T_88294 | conflictPReg_0_12; // @[LoadQueue.scala 192:43:@37807.4]
  assign _T_88296 = _T_88295 | conflictPReg_0_13; // @[LoadQueue.scala 192:43:@37808.4]
  assign _T_88297 = _T_88296 | conflictPReg_0_14; // @[LoadQueue.scala 192:43:@37809.4]
  assign _T_88298 = _T_88297 | conflictPReg_0_15; // @[LoadQueue.scala 192:43:@37810.4]
  assign _GEN_864 = 4'h0 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_865 = 4'h1 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_866 = 4'h2 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_867 = 4'h3 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_868 = 4'h4 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_869 = 4'h5 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_870 = 4'h6 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_871 = 4'h7 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_872 = 4'h8 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_873 = 4'h9 == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_874 = 4'ha == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_875 = 4'hb == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_876 = 4'hc == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_877 = 4'hd == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_878 = 4'he == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_879 = 4'hf == _T_88281; // @[LoadQueue.scala 193:43:@37812.6]
  assign _GEN_881 = 4'h1 == _T_88281 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_882 = 4'h2 == _T_88281 ? shiftedStoreDataKnownPReg_2 : _GEN_881; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_883 = 4'h3 == _T_88281 ? shiftedStoreDataKnownPReg_3 : _GEN_882; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_884 = 4'h4 == _T_88281 ? shiftedStoreDataKnownPReg_4 : _GEN_883; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_885 = 4'h5 == _T_88281 ? shiftedStoreDataKnownPReg_5 : _GEN_884; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_886 = 4'h6 == _T_88281 ? shiftedStoreDataKnownPReg_6 : _GEN_885; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_887 = 4'h7 == _T_88281 ? shiftedStoreDataKnownPReg_7 : _GEN_886; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_888 = 4'h8 == _T_88281 ? shiftedStoreDataKnownPReg_8 : _GEN_887; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_889 = 4'h9 == _T_88281 ? shiftedStoreDataKnownPReg_9 : _GEN_888; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_890 = 4'ha == _T_88281 ? shiftedStoreDataKnownPReg_10 : _GEN_889; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_891 = 4'hb == _T_88281 ? shiftedStoreDataKnownPReg_11 : _GEN_890; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_892 = 4'hc == _T_88281 ? shiftedStoreDataKnownPReg_12 : _GEN_891; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_893 = 4'hd == _T_88281 ? shiftedStoreDataKnownPReg_13 : _GEN_892; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_894 = 4'he == _T_88281 ? shiftedStoreDataKnownPReg_14 : _GEN_893; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_895 = 4'hf == _T_88281 ? shiftedStoreDataKnownPReg_15 : _GEN_894; // @[LoadQueue.scala 194:31:@37813.6]
  assign _GEN_897 = 4'h1 == _T_88281 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_898 = 4'h2 == _T_88281 ? shiftedStoreDataQPreg_2 : _GEN_897; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_899 = 4'h3 == _T_88281 ? shiftedStoreDataQPreg_3 : _GEN_898; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_900 = 4'h4 == _T_88281 ? shiftedStoreDataQPreg_4 : _GEN_899; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_901 = 4'h5 == _T_88281 ? shiftedStoreDataQPreg_5 : _GEN_900; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_902 = 4'h6 == _T_88281 ? shiftedStoreDataQPreg_6 : _GEN_901; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_903 = 4'h7 == _T_88281 ? shiftedStoreDataQPreg_7 : _GEN_902; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_904 = 4'h8 == _T_88281 ? shiftedStoreDataQPreg_8 : _GEN_903; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_905 = 4'h9 == _T_88281 ? shiftedStoreDataQPreg_9 : _GEN_904; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_906 = 4'ha == _T_88281 ? shiftedStoreDataQPreg_10 : _GEN_905; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_907 = 4'hb == _T_88281 ? shiftedStoreDataQPreg_11 : _GEN_906; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_908 = 4'hc == _T_88281 ? shiftedStoreDataQPreg_12 : _GEN_907; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_909 = 4'hd == _T_88281 ? shiftedStoreDataQPreg_13 : _GEN_908; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_910 = 4'he == _T_88281 ? shiftedStoreDataQPreg_14 : _GEN_909; // @[LoadQueue.scala 195:31:@37814.6]
  assign _GEN_911 = 4'hf == _T_88281 ? shiftedStoreDataQPreg_15 : _GEN_910; // @[LoadQueue.scala 195:31:@37814.6]
  assign lastConflict_0_0 = _T_88298 ? _GEN_864 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_1 = _T_88298 ? _GEN_865 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_2 = _T_88298 ? _GEN_866 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_3 = _T_88298 ? _GEN_867 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_4 = _T_88298 ? _GEN_868 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_5 = _T_88298 ? _GEN_869 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_6 = _T_88298 ? _GEN_870 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_7 = _T_88298 ? _GEN_871 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_8 = _T_88298 ? _GEN_872 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_9 = _T_88298 ? _GEN_873 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_10 = _T_88298 ? _GEN_874 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_11 = _T_88298 ? _GEN_875 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_12 = _T_88298 ? _GEN_876 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_13 = _T_88298 ? _GEN_877 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_14 = _T_88298 ? _GEN_878 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign lastConflict_0_15 = _T_88298 ? _GEN_879 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign canBypass_0 = _T_88298 ? _GEN_895 : 1'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign bypassVal_0 = _T_88298 ? _GEN_911 : 32'h0; // @[LoadQueue.scala 192:53:@37811.4]
  assign _T_88404 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[LoadQueue.scala 191:60:@37868.4]
  assign _T_88405 = conflictPReg_1_3 ? 2'h3 : _T_88404; // @[LoadQueue.scala 191:60:@37869.4]
  assign _T_88406 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_88405}; // @[LoadQueue.scala 191:60:@37870.4]
  assign _T_88407 = conflictPReg_1_5 ? 3'h5 : _T_88406; // @[LoadQueue.scala 191:60:@37871.4]
  assign _T_88408 = conflictPReg_1_6 ? 3'h6 : _T_88407; // @[LoadQueue.scala 191:60:@37872.4]
  assign _T_88409 = conflictPReg_1_7 ? 3'h7 : _T_88408; // @[LoadQueue.scala 191:60:@37873.4]
  assign _T_88410 = conflictPReg_1_8 ? 4'h8 : {{1'd0}, _T_88409}; // @[LoadQueue.scala 191:60:@37874.4]
  assign _T_88411 = conflictPReg_1_9 ? 4'h9 : _T_88410; // @[LoadQueue.scala 191:60:@37875.4]
  assign _T_88412 = conflictPReg_1_10 ? 4'ha : _T_88411; // @[LoadQueue.scala 191:60:@37876.4]
  assign _T_88413 = conflictPReg_1_11 ? 4'hb : _T_88412; // @[LoadQueue.scala 191:60:@37877.4]
  assign _T_88414 = conflictPReg_1_12 ? 4'hc : _T_88413; // @[LoadQueue.scala 191:60:@37878.4]
  assign _T_88415 = conflictPReg_1_13 ? 4'hd : _T_88414; // @[LoadQueue.scala 191:60:@37879.4]
  assign _T_88416 = conflictPReg_1_14 ? 4'he : _T_88415; // @[LoadQueue.scala 191:60:@37880.4]
  assign _T_88417 = conflictPReg_1_15 ? 4'hf : _T_88416; // @[LoadQueue.scala 191:60:@37881.4]
  assign _T_88420 = conflictPReg_1_0 | conflictPReg_1_1; // @[LoadQueue.scala 192:43:@37883.4]
  assign _T_88421 = _T_88420 | conflictPReg_1_2; // @[LoadQueue.scala 192:43:@37884.4]
  assign _T_88422 = _T_88421 | conflictPReg_1_3; // @[LoadQueue.scala 192:43:@37885.4]
  assign _T_88423 = _T_88422 | conflictPReg_1_4; // @[LoadQueue.scala 192:43:@37886.4]
  assign _T_88424 = _T_88423 | conflictPReg_1_5; // @[LoadQueue.scala 192:43:@37887.4]
  assign _T_88425 = _T_88424 | conflictPReg_1_6; // @[LoadQueue.scala 192:43:@37888.4]
  assign _T_88426 = _T_88425 | conflictPReg_1_7; // @[LoadQueue.scala 192:43:@37889.4]
  assign _T_88427 = _T_88426 | conflictPReg_1_8; // @[LoadQueue.scala 192:43:@37890.4]
  assign _T_88428 = _T_88427 | conflictPReg_1_9; // @[LoadQueue.scala 192:43:@37891.4]
  assign _T_88429 = _T_88428 | conflictPReg_1_10; // @[LoadQueue.scala 192:43:@37892.4]
  assign _T_88430 = _T_88429 | conflictPReg_1_11; // @[LoadQueue.scala 192:43:@37893.4]
  assign _T_88431 = _T_88430 | conflictPReg_1_12; // @[LoadQueue.scala 192:43:@37894.4]
  assign _T_88432 = _T_88431 | conflictPReg_1_13; // @[LoadQueue.scala 192:43:@37895.4]
  assign _T_88433 = _T_88432 | conflictPReg_1_14; // @[LoadQueue.scala 192:43:@37896.4]
  assign _T_88434 = _T_88433 | conflictPReg_1_15; // @[LoadQueue.scala 192:43:@37897.4]
  assign _GEN_930 = 4'h0 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_931 = 4'h1 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_932 = 4'h2 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_933 = 4'h3 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_934 = 4'h4 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_935 = 4'h5 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_936 = 4'h6 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_937 = 4'h7 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_938 = 4'h8 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_939 = 4'h9 == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_940 = 4'ha == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_941 = 4'hb == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_942 = 4'hc == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_943 = 4'hd == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_944 = 4'he == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_945 = 4'hf == _T_88417; // @[LoadQueue.scala 193:43:@37899.6]
  assign _GEN_947 = 4'h1 == _T_88417 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_948 = 4'h2 == _T_88417 ? shiftedStoreDataKnownPReg_2 : _GEN_947; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_949 = 4'h3 == _T_88417 ? shiftedStoreDataKnownPReg_3 : _GEN_948; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_950 = 4'h4 == _T_88417 ? shiftedStoreDataKnownPReg_4 : _GEN_949; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_951 = 4'h5 == _T_88417 ? shiftedStoreDataKnownPReg_5 : _GEN_950; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_952 = 4'h6 == _T_88417 ? shiftedStoreDataKnownPReg_6 : _GEN_951; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_953 = 4'h7 == _T_88417 ? shiftedStoreDataKnownPReg_7 : _GEN_952; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_954 = 4'h8 == _T_88417 ? shiftedStoreDataKnownPReg_8 : _GEN_953; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_955 = 4'h9 == _T_88417 ? shiftedStoreDataKnownPReg_9 : _GEN_954; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_956 = 4'ha == _T_88417 ? shiftedStoreDataKnownPReg_10 : _GEN_955; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_957 = 4'hb == _T_88417 ? shiftedStoreDataKnownPReg_11 : _GEN_956; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_958 = 4'hc == _T_88417 ? shiftedStoreDataKnownPReg_12 : _GEN_957; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_959 = 4'hd == _T_88417 ? shiftedStoreDataKnownPReg_13 : _GEN_958; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_960 = 4'he == _T_88417 ? shiftedStoreDataKnownPReg_14 : _GEN_959; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_961 = 4'hf == _T_88417 ? shiftedStoreDataKnownPReg_15 : _GEN_960; // @[LoadQueue.scala 194:31:@37900.6]
  assign _GEN_963 = 4'h1 == _T_88417 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_964 = 4'h2 == _T_88417 ? shiftedStoreDataQPreg_2 : _GEN_963; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_965 = 4'h3 == _T_88417 ? shiftedStoreDataQPreg_3 : _GEN_964; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_966 = 4'h4 == _T_88417 ? shiftedStoreDataQPreg_4 : _GEN_965; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_967 = 4'h5 == _T_88417 ? shiftedStoreDataQPreg_5 : _GEN_966; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_968 = 4'h6 == _T_88417 ? shiftedStoreDataQPreg_6 : _GEN_967; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_969 = 4'h7 == _T_88417 ? shiftedStoreDataQPreg_7 : _GEN_968; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_970 = 4'h8 == _T_88417 ? shiftedStoreDataQPreg_8 : _GEN_969; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_971 = 4'h9 == _T_88417 ? shiftedStoreDataQPreg_9 : _GEN_970; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_972 = 4'ha == _T_88417 ? shiftedStoreDataQPreg_10 : _GEN_971; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_973 = 4'hb == _T_88417 ? shiftedStoreDataQPreg_11 : _GEN_972; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_974 = 4'hc == _T_88417 ? shiftedStoreDataQPreg_12 : _GEN_973; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_975 = 4'hd == _T_88417 ? shiftedStoreDataQPreg_13 : _GEN_974; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_976 = 4'he == _T_88417 ? shiftedStoreDataQPreg_14 : _GEN_975; // @[LoadQueue.scala 195:31:@37901.6]
  assign _GEN_977 = 4'hf == _T_88417 ? shiftedStoreDataQPreg_15 : _GEN_976; // @[LoadQueue.scala 195:31:@37901.6]
  assign lastConflict_1_0 = _T_88434 ? _GEN_930 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_1 = _T_88434 ? _GEN_931 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_2 = _T_88434 ? _GEN_932 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_3 = _T_88434 ? _GEN_933 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_4 = _T_88434 ? _GEN_934 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_5 = _T_88434 ? _GEN_935 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_6 = _T_88434 ? _GEN_936 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_7 = _T_88434 ? _GEN_937 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_8 = _T_88434 ? _GEN_938 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_9 = _T_88434 ? _GEN_939 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_10 = _T_88434 ? _GEN_940 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_11 = _T_88434 ? _GEN_941 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_12 = _T_88434 ? _GEN_942 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_13 = _T_88434 ? _GEN_943 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_14 = _T_88434 ? _GEN_944 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign lastConflict_1_15 = _T_88434 ? _GEN_945 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign canBypass_1 = _T_88434 ? _GEN_961 : 1'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign bypassVal_1 = _T_88434 ? _GEN_977 : 32'h0; // @[LoadQueue.scala 192:53:@37898.4]
  assign _T_88540 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[LoadQueue.scala 191:60:@37955.4]
  assign _T_88541 = conflictPReg_2_3 ? 2'h3 : _T_88540; // @[LoadQueue.scala 191:60:@37956.4]
  assign _T_88542 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_88541}; // @[LoadQueue.scala 191:60:@37957.4]
  assign _T_88543 = conflictPReg_2_5 ? 3'h5 : _T_88542; // @[LoadQueue.scala 191:60:@37958.4]
  assign _T_88544 = conflictPReg_2_6 ? 3'h6 : _T_88543; // @[LoadQueue.scala 191:60:@37959.4]
  assign _T_88545 = conflictPReg_2_7 ? 3'h7 : _T_88544; // @[LoadQueue.scala 191:60:@37960.4]
  assign _T_88546 = conflictPReg_2_8 ? 4'h8 : {{1'd0}, _T_88545}; // @[LoadQueue.scala 191:60:@37961.4]
  assign _T_88547 = conflictPReg_2_9 ? 4'h9 : _T_88546; // @[LoadQueue.scala 191:60:@37962.4]
  assign _T_88548 = conflictPReg_2_10 ? 4'ha : _T_88547; // @[LoadQueue.scala 191:60:@37963.4]
  assign _T_88549 = conflictPReg_2_11 ? 4'hb : _T_88548; // @[LoadQueue.scala 191:60:@37964.4]
  assign _T_88550 = conflictPReg_2_12 ? 4'hc : _T_88549; // @[LoadQueue.scala 191:60:@37965.4]
  assign _T_88551 = conflictPReg_2_13 ? 4'hd : _T_88550; // @[LoadQueue.scala 191:60:@37966.4]
  assign _T_88552 = conflictPReg_2_14 ? 4'he : _T_88551; // @[LoadQueue.scala 191:60:@37967.4]
  assign _T_88553 = conflictPReg_2_15 ? 4'hf : _T_88552; // @[LoadQueue.scala 191:60:@37968.4]
  assign _T_88556 = conflictPReg_2_0 | conflictPReg_2_1; // @[LoadQueue.scala 192:43:@37970.4]
  assign _T_88557 = _T_88556 | conflictPReg_2_2; // @[LoadQueue.scala 192:43:@37971.4]
  assign _T_88558 = _T_88557 | conflictPReg_2_3; // @[LoadQueue.scala 192:43:@37972.4]
  assign _T_88559 = _T_88558 | conflictPReg_2_4; // @[LoadQueue.scala 192:43:@37973.4]
  assign _T_88560 = _T_88559 | conflictPReg_2_5; // @[LoadQueue.scala 192:43:@37974.4]
  assign _T_88561 = _T_88560 | conflictPReg_2_6; // @[LoadQueue.scala 192:43:@37975.4]
  assign _T_88562 = _T_88561 | conflictPReg_2_7; // @[LoadQueue.scala 192:43:@37976.4]
  assign _T_88563 = _T_88562 | conflictPReg_2_8; // @[LoadQueue.scala 192:43:@37977.4]
  assign _T_88564 = _T_88563 | conflictPReg_2_9; // @[LoadQueue.scala 192:43:@37978.4]
  assign _T_88565 = _T_88564 | conflictPReg_2_10; // @[LoadQueue.scala 192:43:@37979.4]
  assign _T_88566 = _T_88565 | conflictPReg_2_11; // @[LoadQueue.scala 192:43:@37980.4]
  assign _T_88567 = _T_88566 | conflictPReg_2_12; // @[LoadQueue.scala 192:43:@37981.4]
  assign _T_88568 = _T_88567 | conflictPReg_2_13; // @[LoadQueue.scala 192:43:@37982.4]
  assign _T_88569 = _T_88568 | conflictPReg_2_14; // @[LoadQueue.scala 192:43:@37983.4]
  assign _T_88570 = _T_88569 | conflictPReg_2_15; // @[LoadQueue.scala 192:43:@37984.4]
  assign _GEN_996 = 4'h0 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_997 = 4'h1 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_998 = 4'h2 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_999 = 4'h3 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1000 = 4'h4 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1001 = 4'h5 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1002 = 4'h6 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1003 = 4'h7 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1004 = 4'h8 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1005 = 4'h9 == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1006 = 4'ha == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1007 = 4'hb == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1008 = 4'hc == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1009 = 4'hd == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1010 = 4'he == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1011 = 4'hf == _T_88553; // @[LoadQueue.scala 193:43:@37986.6]
  assign _GEN_1013 = 4'h1 == _T_88553 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1014 = 4'h2 == _T_88553 ? shiftedStoreDataKnownPReg_2 : _GEN_1013; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1015 = 4'h3 == _T_88553 ? shiftedStoreDataKnownPReg_3 : _GEN_1014; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1016 = 4'h4 == _T_88553 ? shiftedStoreDataKnownPReg_4 : _GEN_1015; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1017 = 4'h5 == _T_88553 ? shiftedStoreDataKnownPReg_5 : _GEN_1016; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1018 = 4'h6 == _T_88553 ? shiftedStoreDataKnownPReg_6 : _GEN_1017; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1019 = 4'h7 == _T_88553 ? shiftedStoreDataKnownPReg_7 : _GEN_1018; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1020 = 4'h8 == _T_88553 ? shiftedStoreDataKnownPReg_8 : _GEN_1019; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1021 = 4'h9 == _T_88553 ? shiftedStoreDataKnownPReg_9 : _GEN_1020; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1022 = 4'ha == _T_88553 ? shiftedStoreDataKnownPReg_10 : _GEN_1021; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1023 = 4'hb == _T_88553 ? shiftedStoreDataKnownPReg_11 : _GEN_1022; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1024 = 4'hc == _T_88553 ? shiftedStoreDataKnownPReg_12 : _GEN_1023; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1025 = 4'hd == _T_88553 ? shiftedStoreDataKnownPReg_13 : _GEN_1024; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1026 = 4'he == _T_88553 ? shiftedStoreDataKnownPReg_14 : _GEN_1025; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1027 = 4'hf == _T_88553 ? shiftedStoreDataKnownPReg_15 : _GEN_1026; // @[LoadQueue.scala 194:31:@37987.6]
  assign _GEN_1029 = 4'h1 == _T_88553 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1030 = 4'h2 == _T_88553 ? shiftedStoreDataQPreg_2 : _GEN_1029; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1031 = 4'h3 == _T_88553 ? shiftedStoreDataQPreg_3 : _GEN_1030; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1032 = 4'h4 == _T_88553 ? shiftedStoreDataQPreg_4 : _GEN_1031; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1033 = 4'h5 == _T_88553 ? shiftedStoreDataQPreg_5 : _GEN_1032; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1034 = 4'h6 == _T_88553 ? shiftedStoreDataQPreg_6 : _GEN_1033; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1035 = 4'h7 == _T_88553 ? shiftedStoreDataQPreg_7 : _GEN_1034; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1036 = 4'h8 == _T_88553 ? shiftedStoreDataQPreg_8 : _GEN_1035; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1037 = 4'h9 == _T_88553 ? shiftedStoreDataQPreg_9 : _GEN_1036; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1038 = 4'ha == _T_88553 ? shiftedStoreDataQPreg_10 : _GEN_1037; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1039 = 4'hb == _T_88553 ? shiftedStoreDataQPreg_11 : _GEN_1038; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1040 = 4'hc == _T_88553 ? shiftedStoreDataQPreg_12 : _GEN_1039; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1041 = 4'hd == _T_88553 ? shiftedStoreDataQPreg_13 : _GEN_1040; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1042 = 4'he == _T_88553 ? shiftedStoreDataQPreg_14 : _GEN_1041; // @[LoadQueue.scala 195:31:@37988.6]
  assign _GEN_1043 = 4'hf == _T_88553 ? shiftedStoreDataQPreg_15 : _GEN_1042; // @[LoadQueue.scala 195:31:@37988.6]
  assign lastConflict_2_0 = _T_88570 ? _GEN_996 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_1 = _T_88570 ? _GEN_997 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_2 = _T_88570 ? _GEN_998 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_3 = _T_88570 ? _GEN_999 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_4 = _T_88570 ? _GEN_1000 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_5 = _T_88570 ? _GEN_1001 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_6 = _T_88570 ? _GEN_1002 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_7 = _T_88570 ? _GEN_1003 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_8 = _T_88570 ? _GEN_1004 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_9 = _T_88570 ? _GEN_1005 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_10 = _T_88570 ? _GEN_1006 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_11 = _T_88570 ? _GEN_1007 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_12 = _T_88570 ? _GEN_1008 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_13 = _T_88570 ? _GEN_1009 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_14 = _T_88570 ? _GEN_1010 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign lastConflict_2_15 = _T_88570 ? _GEN_1011 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign canBypass_2 = _T_88570 ? _GEN_1027 : 1'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign bypassVal_2 = _T_88570 ? _GEN_1043 : 32'h0; // @[LoadQueue.scala 192:53:@37985.4]
  assign _T_88676 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[LoadQueue.scala 191:60:@38042.4]
  assign _T_88677 = conflictPReg_3_3 ? 2'h3 : _T_88676; // @[LoadQueue.scala 191:60:@38043.4]
  assign _T_88678 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_88677}; // @[LoadQueue.scala 191:60:@38044.4]
  assign _T_88679 = conflictPReg_3_5 ? 3'h5 : _T_88678; // @[LoadQueue.scala 191:60:@38045.4]
  assign _T_88680 = conflictPReg_3_6 ? 3'h6 : _T_88679; // @[LoadQueue.scala 191:60:@38046.4]
  assign _T_88681 = conflictPReg_3_7 ? 3'h7 : _T_88680; // @[LoadQueue.scala 191:60:@38047.4]
  assign _T_88682 = conflictPReg_3_8 ? 4'h8 : {{1'd0}, _T_88681}; // @[LoadQueue.scala 191:60:@38048.4]
  assign _T_88683 = conflictPReg_3_9 ? 4'h9 : _T_88682; // @[LoadQueue.scala 191:60:@38049.4]
  assign _T_88684 = conflictPReg_3_10 ? 4'ha : _T_88683; // @[LoadQueue.scala 191:60:@38050.4]
  assign _T_88685 = conflictPReg_3_11 ? 4'hb : _T_88684; // @[LoadQueue.scala 191:60:@38051.4]
  assign _T_88686 = conflictPReg_3_12 ? 4'hc : _T_88685; // @[LoadQueue.scala 191:60:@38052.4]
  assign _T_88687 = conflictPReg_3_13 ? 4'hd : _T_88686; // @[LoadQueue.scala 191:60:@38053.4]
  assign _T_88688 = conflictPReg_3_14 ? 4'he : _T_88687; // @[LoadQueue.scala 191:60:@38054.4]
  assign _T_88689 = conflictPReg_3_15 ? 4'hf : _T_88688; // @[LoadQueue.scala 191:60:@38055.4]
  assign _T_88692 = conflictPReg_3_0 | conflictPReg_3_1; // @[LoadQueue.scala 192:43:@38057.4]
  assign _T_88693 = _T_88692 | conflictPReg_3_2; // @[LoadQueue.scala 192:43:@38058.4]
  assign _T_88694 = _T_88693 | conflictPReg_3_3; // @[LoadQueue.scala 192:43:@38059.4]
  assign _T_88695 = _T_88694 | conflictPReg_3_4; // @[LoadQueue.scala 192:43:@38060.4]
  assign _T_88696 = _T_88695 | conflictPReg_3_5; // @[LoadQueue.scala 192:43:@38061.4]
  assign _T_88697 = _T_88696 | conflictPReg_3_6; // @[LoadQueue.scala 192:43:@38062.4]
  assign _T_88698 = _T_88697 | conflictPReg_3_7; // @[LoadQueue.scala 192:43:@38063.4]
  assign _T_88699 = _T_88698 | conflictPReg_3_8; // @[LoadQueue.scala 192:43:@38064.4]
  assign _T_88700 = _T_88699 | conflictPReg_3_9; // @[LoadQueue.scala 192:43:@38065.4]
  assign _T_88701 = _T_88700 | conflictPReg_3_10; // @[LoadQueue.scala 192:43:@38066.4]
  assign _T_88702 = _T_88701 | conflictPReg_3_11; // @[LoadQueue.scala 192:43:@38067.4]
  assign _T_88703 = _T_88702 | conflictPReg_3_12; // @[LoadQueue.scala 192:43:@38068.4]
  assign _T_88704 = _T_88703 | conflictPReg_3_13; // @[LoadQueue.scala 192:43:@38069.4]
  assign _T_88705 = _T_88704 | conflictPReg_3_14; // @[LoadQueue.scala 192:43:@38070.4]
  assign _T_88706 = _T_88705 | conflictPReg_3_15; // @[LoadQueue.scala 192:43:@38071.4]
  assign _GEN_1062 = 4'h0 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1063 = 4'h1 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1064 = 4'h2 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1065 = 4'h3 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1066 = 4'h4 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1067 = 4'h5 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1068 = 4'h6 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1069 = 4'h7 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1070 = 4'h8 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1071 = 4'h9 == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1072 = 4'ha == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1073 = 4'hb == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1074 = 4'hc == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1075 = 4'hd == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1076 = 4'he == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1077 = 4'hf == _T_88689; // @[LoadQueue.scala 193:43:@38073.6]
  assign _GEN_1079 = 4'h1 == _T_88689 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1080 = 4'h2 == _T_88689 ? shiftedStoreDataKnownPReg_2 : _GEN_1079; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1081 = 4'h3 == _T_88689 ? shiftedStoreDataKnownPReg_3 : _GEN_1080; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1082 = 4'h4 == _T_88689 ? shiftedStoreDataKnownPReg_4 : _GEN_1081; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1083 = 4'h5 == _T_88689 ? shiftedStoreDataKnownPReg_5 : _GEN_1082; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1084 = 4'h6 == _T_88689 ? shiftedStoreDataKnownPReg_6 : _GEN_1083; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1085 = 4'h7 == _T_88689 ? shiftedStoreDataKnownPReg_7 : _GEN_1084; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1086 = 4'h8 == _T_88689 ? shiftedStoreDataKnownPReg_8 : _GEN_1085; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1087 = 4'h9 == _T_88689 ? shiftedStoreDataKnownPReg_9 : _GEN_1086; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1088 = 4'ha == _T_88689 ? shiftedStoreDataKnownPReg_10 : _GEN_1087; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1089 = 4'hb == _T_88689 ? shiftedStoreDataKnownPReg_11 : _GEN_1088; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1090 = 4'hc == _T_88689 ? shiftedStoreDataKnownPReg_12 : _GEN_1089; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1091 = 4'hd == _T_88689 ? shiftedStoreDataKnownPReg_13 : _GEN_1090; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1092 = 4'he == _T_88689 ? shiftedStoreDataKnownPReg_14 : _GEN_1091; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1093 = 4'hf == _T_88689 ? shiftedStoreDataKnownPReg_15 : _GEN_1092; // @[LoadQueue.scala 194:31:@38074.6]
  assign _GEN_1095 = 4'h1 == _T_88689 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1096 = 4'h2 == _T_88689 ? shiftedStoreDataQPreg_2 : _GEN_1095; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1097 = 4'h3 == _T_88689 ? shiftedStoreDataQPreg_3 : _GEN_1096; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1098 = 4'h4 == _T_88689 ? shiftedStoreDataQPreg_4 : _GEN_1097; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1099 = 4'h5 == _T_88689 ? shiftedStoreDataQPreg_5 : _GEN_1098; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1100 = 4'h6 == _T_88689 ? shiftedStoreDataQPreg_6 : _GEN_1099; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1101 = 4'h7 == _T_88689 ? shiftedStoreDataQPreg_7 : _GEN_1100; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1102 = 4'h8 == _T_88689 ? shiftedStoreDataQPreg_8 : _GEN_1101; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1103 = 4'h9 == _T_88689 ? shiftedStoreDataQPreg_9 : _GEN_1102; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1104 = 4'ha == _T_88689 ? shiftedStoreDataQPreg_10 : _GEN_1103; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1105 = 4'hb == _T_88689 ? shiftedStoreDataQPreg_11 : _GEN_1104; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1106 = 4'hc == _T_88689 ? shiftedStoreDataQPreg_12 : _GEN_1105; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1107 = 4'hd == _T_88689 ? shiftedStoreDataQPreg_13 : _GEN_1106; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1108 = 4'he == _T_88689 ? shiftedStoreDataQPreg_14 : _GEN_1107; // @[LoadQueue.scala 195:31:@38075.6]
  assign _GEN_1109 = 4'hf == _T_88689 ? shiftedStoreDataQPreg_15 : _GEN_1108; // @[LoadQueue.scala 195:31:@38075.6]
  assign lastConflict_3_0 = _T_88706 ? _GEN_1062 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_1 = _T_88706 ? _GEN_1063 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_2 = _T_88706 ? _GEN_1064 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_3 = _T_88706 ? _GEN_1065 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_4 = _T_88706 ? _GEN_1066 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_5 = _T_88706 ? _GEN_1067 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_6 = _T_88706 ? _GEN_1068 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_7 = _T_88706 ? _GEN_1069 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_8 = _T_88706 ? _GEN_1070 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_9 = _T_88706 ? _GEN_1071 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_10 = _T_88706 ? _GEN_1072 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_11 = _T_88706 ? _GEN_1073 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_12 = _T_88706 ? _GEN_1074 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_13 = _T_88706 ? _GEN_1075 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_14 = _T_88706 ? _GEN_1076 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign lastConflict_3_15 = _T_88706 ? _GEN_1077 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign canBypass_3 = _T_88706 ? _GEN_1093 : 1'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign bypassVal_3 = _T_88706 ? _GEN_1109 : 32'h0; // @[LoadQueue.scala 192:53:@38072.4]
  assign _T_88812 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[LoadQueue.scala 191:60:@38129.4]
  assign _T_88813 = conflictPReg_4_3 ? 2'h3 : _T_88812; // @[LoadQueue.scala 191:60:@38130.4]
  assign _T_88814 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_88813}; // @[LoadQueue.scala 191:60:@38131.4]
  assign _T_88815 = conflictPReg_4_5 ? 3'h5 : _T_88814; // @[LoadQueue.scala 191:60:@38132.4]
  assign _T_88816 = conflictPReg_4_6 ? 3'h6 : _T_88815; // @[LoadQueue.scala 191:60:@38133.4]
  assign _T_88817 = conflictPReg_4_7 ? 3'h7 : _T_88816; // @[LoadQueue.scala 191:60:@38134.4]
  assign _T_88818 = conflictPReg_4_8 ? 4'h8 : {{1'd0}, _T_88817}; // @[LoadQueue.scala 191:60:@38135.4]
  assign _T_88819 = conflictPReg_4_9 ? 4'h9 : _T_88818; // @[LoadQueue.scala 191:60:@38136.4]
  assign _T_88820 = conflictPReg_4_10 ? 4'ha : _T_88819; // @[LoadQueue.scala 191:60:@38137.4]
  assign _T_88821 = conflictPReg_4_11 ? 4'hb : _T_88820; // @[LoadQueue.scala 191:60:@38138.4]
  assign _T_88822 = conflictPReg_4_12 ? 4'hc : _T_88821; // @[LoadQueue.scala 191:60:@38139.4]
  assign _T_88823 = conflictPReg_4_13 ? 4'hd : _T_88822; // @[LoadQueue.scala 191:60:@38140.4]
  assign _T_88824 = conflictPReg_4_14 ? 4'he : _T_88823; // @[LoadQueue.scala 191:60:@38141.4]
  assign _T_88825 = conflictPReg_4_15 ? 4'hf : _T_88824; // @[LoadQueue.scala 191:60:@38142.4]
  assign _T_88828 = conflictPReg_4_0 | conflictPReg_4_1; // @[LoadQueue.scala 192:43:@38144.4]
  assign _T_88829 = _T_88828 | conflictPReg_4_2; // @[LoadQueue.scala 192:43:@38145.4]
  assign _T_88830 = _T_88829 | conflictPReg_4_3; // @[LoadQueue.scala 192:43:@38146.4]
  assign _T_88831 = _T_88830 | conflictPReg_4_4; // @[LoadQueue.scala 192:43:@38147.4]
  assign _T_88832 = _T_88831 | conflictPReg_4_5; // @[LoadQueue.scala 192:43:@38148.4]
  assign _T_88833 = _T_88832 | conflictPReg_4_6; // @[LoadQueue.scala 192:43:@38149.4]
  assign _T_88834 = _T_88833 | conflictPReg_4_7; // @[LoadQueue.scala 192:43:@38150.4]
  assign _T_88835 = _T_88834 | conflictPReg_4_8; // @[LoadQueue.scala 192:43:@38151.4]
  assign _T_88836 = _T_88835 | conflictPReg_4_9; // @[LoadQueue.scala 192:43:@38152.4]
  assign _T_88837 = _T_88836 | conflictPReg_4_10; // @[LoadQueue.scala 192:43:@38153.4]
  assign _T_88838 = _T_88837 | conflictPReg_4_11; // @[LoadQueue.scala 192:43:@38154.4]
  assign _T_88839 = _T_88838 | conflictPReg_4_12; // @[LoadQueue.scala 192:43:@38155.4]
  assign _T_88840 = _T_88839 | conflictPReg_4_13; // @[LoadQueue.scala 192:43:@38156.4]
  assign _T_88841 = _T_88840 | conflictPReg_4_14; // @[LoadQueue.scala 192:43:@38157.4]
  assign _T_88842 = _T_88841 | conflictPReg_4_15; // @[LoadQueue.scala 192:43:@38158.4]
  assign _GEN_1128 = 4'h0 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1129 = 4'h1 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1130 = 4'h2 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1131 = 4'h3 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1132 = 4'h4 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1133 = 4'h5 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1134 = 4'h6 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1135 = 4'h7 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1136 = 4'h8 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1137 = 4'h9 == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1138 = 4'ha == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1139 = 4'hb == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1140 = 4'hc == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1141 = 4'hd == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1142 = 4'he == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1143 = 4'hf == _T_88825; // @[LoadQueue.scala 193:43:@38160.6]
  assign _GEN_1145 = 4'h1 == _T_88825 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1146 = 4'h2 == _T_88825 ? shiftedStoreDataKnownPReg_2 : _GEN_1145; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1147 = 4'h3 == _T_88825 ? shiftedStoreDataKnownPReg_3 : _GEN_1146; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1148 = 4'h4 == _T_88825 ? shiftedStoreDataKnownPReg_4 : _GEN_1147; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1149 = 4'h5 == _T_88825 ? shiftedStoreDataKnownPReg_5 : _GEN_1148; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1150 = 4'h6 == _T_88825 ? shiftedStoreDataKnownPReg_6 : _GEN_1149; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1151 = 4'h7 == _T_88825 ? shiftedStoreDataKnownPReg_7 : _GEN_1150; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1152 = 4'h8 == _T_88825 ? shiftedStoreDataKnownPReg_8 : _GEN_1151; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1153 = 4'h9 == _T_88825 ? shiftedStoreDataKnownPReg_9 : _GEN_1152; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1154 = 4'ha == _T_88825 ? shiftedStoreDataKnownPReg_10 : _GEN_1153; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1155 = 4'hb == _T_88825 ? shiftedStoreDataKnownPReg_11 : _GEN_1154; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1156 = 4'hc == _T_88825 ? shiftedStoreDataKnownPReg_12 : _GEN_1155; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1157 = 4'hd == _T_88825 ? shiftedStoreDataKnownPReg_13 : _GEN_1156; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1158 = 4'he == _T_88825 ? shiftedStoreDataKnownPReg_14 : _GEN_1157; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1159 = 4'hf == _T_88825 ? shiftedStoreDataKnownPReg_15 : _GEN_1158; // @[LoadQueue.scala 194:31:@38161.6]
  assign _GEN_1161 = 4'h1 == _T_88825 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1162 = 4'h2 == _T_88825 ? shiftedStoreDataQPreg_2 : _GEN_1161; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1163 = 4'h3 == _T_88825 ? shiftedStoreDataQPreg_3 : _GEN_1162; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1164 = 4'h4 == _T_88825 ? shiftedStoreDataQPreg_4 : _GEN_1163; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1165 = 4'h5 == _T_88825 ? shiftedStoreDataQPreg_5 : _GEN_1164; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1166 = 4'h6 == _T_88825 ? shiftedStoreDataQPreg_6 : _GEN_1165; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1167 = 4'h7 == _T_88825 ? shiftedStoreDataQPreg_7 : _GEN_1166; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1168 = 4'h8 == _T_88825 ? shiftedStoreDataQPreg_8 : _GEN_1167; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1169 = 4'h9 == _T_88825 ? shiftedStoreDataQPreg_9 : _GEN_1168; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1170 = 4'ha == _T_88825 ? shiftedStoreDataQPreg_10 : _GEN_1169; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1171 = 4'hb == _T_88825 ? shiftedStoreDataQPreg_11 : _GEN_1170; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1172 = 4'hc == _T_88825 ? shiftedStoreDataQPreg_12 : _GEN_1171; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1173 = 4'hd == _T_88825 ? shiftedStoreDataQPreg_13 : _GEN_1172; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1174 = 4'he == _T_88825 ? shiftedStoreDataQPreg_14 : _GEN_1173; // @[LoadQueue.scala 195:31:@38162.6]
  assign _GEN_1175 = 4'hf == _T_88825 ? shiftedStoreDataQPreg_15 : _GEN_1174; // @[LoadQueue.scala 195:31:@38162.6]
  assign lastConflict_4_0 = _T_88842 ? _GEN_1128 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_1 = _T_88842 ? _GEN_1129 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_2 = _T_88842 ? _GEN_1130 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_3 = _T_88842 ? _GEN_1131 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_4 = _T_88842 ? _GEN_1132 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_5 = _T_88842 ? _GEN_1133 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_6 = _T_88842 ? _GEN_1134 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_7 = _T_88842 ? _GEN_1135 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_8 = _T_88842 ? _GEN_1136 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_9 = _T_88842 ? _GEN_1137 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_10 = _T_88842 ? _GEN_1138 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_11 = _T_88842 ? _GEN_1139 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_12 = _T_88842 ? _GEN_1140 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_13 = _T_88842 ? _GEN_1141 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_14 = _T_88842 ? _GEN_1142 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign lastConflict_4_15 = _T_88842 ? _GEN_1143 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign canBypass_4 = _T_88842 ? _GEN_1159 : 1'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign bypassVal_4 = _T_88842 ? _GEN_1175 : 32'h0; // @[LoadQueue.scala 192:53:@38159.4]
  assign _T_88948 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[LoadQueue.scala 191:60:@38216.4]
  assign _T_88949 = conflictPReg_5_3 ? 2'h3 : _T_88948; // @[LoadQueue.scala 191:60:@38217.4]
  assign _T_88950 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_88949}; // @[LoadQueue.scala 191:60:@38218.4]
  assign _T_88951 = conflictPReg_5_5 ? 3'h5 : _T_88950; // @[LoadQueue.scala 191:60:@38219.4]
  assign _T_88952 = conflictPReg_5_6 ? 3'h6 : _T_88951; // @[LoadQueue.scala 191:60:@38220.4]
  assign _T_88953 = conflictPReg_5_7 ? 3'h7 : _T_88952; // @[LoadQueue.scala 191:60:@38221.4]
  assign _T_88954 = conflictPReg_5_8 ? 4'h8 : {{1'd0}, _T_88953}; // @[LoadQueue.scala 191:60:@38222.4]
  assign _T_88955 = conflictPReg_5_9 ? 4'h9 : _T_88954; // @[LoadQueue.scala 191:60:@38223.4]
  assign _T_88956 = conflictPReg_5_10 ? 4'ha : _T_88955; // @[LoadQueue.scala 191:60:@38224.4]
  assign _T_88957 = conflictPReg_5_11 ? 4'hb : _T_88956; // @[LoadQueue.scala 191:60:@38225.4]
  assign _T_88958 = conflictPReg_5_12 ? 4'hc : _T_88957; // @[LoadQueue.scala 191:60:@38226.4]
  assign _T_88959 = conflictPReg_5_13 ? 4'hd : _T_88958; // @[LoadQueue.scala 191:60:@38227.4]
  assign _T_88960 = conflictPReg_5_14 ? 4'he : _T_88959; // @[LoadQueue.scala 191:60:@38228.4]
  assign _T_88961 = conflictPReg_5_15 ? 4'hf : _T_88960; // @[LoadQueue.scala 191:60:@38229.4]
  assign _T_88964 = conflictPReg_5_0 | conflictPReg_5_1; // @[LoadQueue.scala 192:43:@38231.4]
  assign _T_88965 = _T_88964 | conflictPReg_5_2; // @[LoadQueue.scala 192:43:@38232.4]
  assign _T_88966 = _T_88965 | conflictPReg_5_3; // @[LoadQueue.scala 192:43:@38233.4]
  assign _T_88967 = _T_88966 | conflictPReg_5_4; // @[LoadQueue.scala 192:43:@38234.4]
  assign _T_88968 = _T_88967 | conflictPReg_5_5; // @[LoadQueue.scala 192:43:@38235.4]
  assign _T_88969 = _T_88968 | conflictPReg_5_6; // @[LoadQueue.scala 192:43:@38236.4]
  assign _T_88970 = _T_88969 | conflictPReg_5_7; // @[LoadQueue.scala 192:43:@38237.4]
  assign _T_88971 = _T_88970 | conflictPReg_5_8; // @[LoadQueue.scala 192:43:@38238.4]
  assign _T_88972 = _T_88971 | conflictPReg_5_9; // @[LoadQueue.scala 192:43:@38239.4]
  assign _T_88973 = _T_88972 | conflictPReg_5_10; // @[LoadQueue.scala 192:43:@38240.4]
  assign _T_88974 = _T_88973 | conflictPReg_5_11; // @[LoadQueue.scala 192:43:@38241.4]
  assign _T_88975 = _T_88974 | conflictPReg_5_12; // @[LoadQueue.scala 192:43:@38242.4]
  assign _T_88976 = _T_88975 | conflictPReg_5_13; // @[LoadQueue.scala 192:43:@38243.4]
  assign _T_88977 = _T_88976 | conflictPReg_5_14; // @[LoadQueue.scala 192:43:@38244.4]
  assign _T_88978 = _T_88977 | conflictPReg_5_15; // @[LoadQueue.scala 192:43:@38245.4]
  assign _GEN_1194 = 4'h0 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1195 = 4'h1 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1196 = 4'h2 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1197 = 4'h3 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1198 = 4'h4 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1199 = 4'h5 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1200 = 4'h6 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1201 = 4'h7 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1202 = 4'h8 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1203 = 4'h9 == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1204 = 4'ha == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1205 = 4'hb == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1206 = 4'hc == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1207 = 4'hd == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1208 = 4'he == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1209 = 4'hf == _T_88961; // @[LoadQueue.scala 193:43:@38247.6]
  assign _GEN_1211 = 4'h1 == _T_88961 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1212 = 4'h2 == _T_88961 ? shiftedStoreDataKnownPReg_2 : _GEN_1211; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1213 = 4'h3 == _T_88961 ? shiftedStoreDataKnownPReg_3 : _GEN_1212; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1214 = 4'h4 == _T_88961 ? shiftedStoreDataKnownPReg_4 : _GEN_1213; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1215 = 4'h5 == _T_88961 ? shiftedStoreDataKnownPReg_5 : _GEN_1214; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1216 = 4'h6 == _T_88961 ? shiftedStoreDataKnownPReg_6 : _GEN_1215; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1217 = 4'h7 == _T_88961 ? shiftedStoreDataKnownPReg_7 : _GEN_1216; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1218 = 4'h8 == _T_88961 ? shiftedStoreDataKnownPReg_8 : _GEN_1217; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1219 = 4'h9 == _T_88961 ? shiftedStoreDataKnownPReg_9 : _GEN_1218; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1220 = 4'ha == _T_88961 ? shiftedStoreDataKnownPReg_10 : _GEN_1219; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1221 = 4'hb == _T_88961 ? shiftedStoreDataKnownPReg_11 : _GEN_1220; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1222 = 4'hc == _T_88961 ? shiftedStoreDataKnownPReg_12 : _GEN_1221; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1223 = 4'hd == _T_88961 ? shiftedStoreDataKnownPReg_13 : _GEN_1222; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1224 = 4'he == _T_88961 ? shiftedStoreDataKnownPReg_14 : _GEN_1223; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1225 = 4'hf == _T_88961 ? shiftedStoreDataKnownPReg_15 : _GEN_1224; // @[LoadQueue.scala 194:31:@38248.6]
  assign _GEN_1227 = 4'h1 == _T_88961 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1228 = 4'h2 == _T_88961 ? shiftedStoreDataQPreg_2 : _GEN_1227; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1229 = 4'h3 == _T_88961 ? shiftedStoreDataQPreg_3 : _GEN_1228; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1230 = 4'h4 == _T_88961 ? shiftedStoreDataQPreg_4 : _GEN_1229; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1231 = 4'h5 == _T_88961 ? shiftedStoreDataQPreg_5 : _GEN_1230; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1232 = 4'h6 == _T_88961 ? shiftedStoreDataQPreg_6 : _GEN_1231; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1233 = 4'h7 == _T_88961 ? shiftedStoreDataQPreg_7 : _GEN_1232; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1234 = 4'h8 == _T_88961 ? shiftedStoreDataQPreg_8 : _GEN_1233; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1235 = 4'h9 == _T_88961 ? shiftedStoreDataQPreg_9 : _GEN_1234; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1236 = 4'ha == _T_88961 ? shiftedStoreDataQPreg_10 : _GEN_1235; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1237 = 4'hb == _T_88961 ? shiftedStoreDataQPreg_11 : _GEN_1236; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1238 = 4'hc == _T_88961 ? shiftedStoreDataQPreg_12 : _GEN_1237; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1239 = 4'hd == _T_88961 ? shiftedStoreDataQPreg_13 : _GEN_1238; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1240 = 4'he == _T_88961 ? shiftedStoreDataQPreg_14 : _GEN_1239; // @[LoadQueue.scala 195:31:@38249.6]
  assign _GEN_1241 = 4'hf == _T_88961 ? shiftedStoreDataQPreg_15 : _GEN_1240; // @[LoadQueue.scala 195:31:@38249.6]
  assign lastConflict_5_0 = _T_88978 ? _GEN_1194 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_1 = _T_88978 ? _GEN_1195 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_2 = _T_88978 ? _GEN_1196 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_3 = _T_88978 ? _GEN_1197 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_4 = _T_88978 ? _GEN_1198 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_5 = _T_88978 ? _GEN_1199 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_6 = _T_88978 ? _GEN_1200 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_7 = _T_88978 ? _GEN_1201 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_8 = _T_88978 ? _GEN_1202 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_9 = _T_88978 ? _GEN_1203 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_10 = _T_88978 ? _GEN_1204 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_11 = _T_88978 ? _GEN_1205 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_12 = _T_88978 ? _GEN_1206 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_13 = _T_88978 ? _GEN_1207 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_14 = _T_88978 ? _GEN_1208 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign lastConflict_5_15 = _T_88978 ? _GEN_1209 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign canBypass_5 = _T_88978 ? _GEN_1225 : 1'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign bypassVal_5 = _T_88978 ? _GEN_1241 : 32'h0; // @[LoadQueue.scala 192:53:@38246.4]
  assign _T_89084 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[LoadQueue.scala 191:60:@38303.4]
  assign _T_89085 = conflictPReg_6_3 ? 2'h3 : _T_89084; // @[LoadQueue.scala 191:60:@38304.4]
  assign _T_89086 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_89085}; // @[LoadQueue.scala 191:60:@38305.4]
  assign _T_89087 = conflictPReg_6_5 ? 3'h5 : _T_89086; // @[LoadQueue.scala 191:60:@38306.4]
  assign _T_89088 = conflictPReg_6_6 ? 3'h6 : _T_89087; // @[LoadQueue.scala 191:60:@38307.4]
  assign _T_89089 = conflictPReg_6_7 ? 3'h7 : _T_89088; // @[LoadQueue.scala 191:60:@38308.4]
  assign _T_89090 = conflictPReg_6_8 ? 4'h8 : {{1'd0}, _T_89089}; // @[LoadQueue.scala 191:60:@38309.4]
  assign _T_89091 = conflictPReg_6_9 ? 4'h9 : _T_89090; // @[LoadQueue.scala 191:60:@38310.4]
  assign _T_89092 = conflictPReg_6_10 ? 4'ha : _T_89091; // @[LoadQueue.scala 191:60:@38311.4]
  assign _T_89093 = conflictPReg_6_11 ? 4'hb : _T_89092; // @[LoadQueue.scala 191:60:@38312.4]
  assign _T_89094 = conflictPReg_6_12 ? 4'hc : _T_89093; // @[LoadQueue.scala 191:60:@38313.4]
  assign _T_89095 = conflictPReg_6_13 ? 4'hd : _T_89094; // @[LoadQueue.scala 191:60:@38314.4]
  assign _T_89096 = conflictPReg_6_14 ? 4'he : _T_89095; // @[LoadQueue.scala 191:60:@38315.4]
  assign _T_89097 = conflictPReg_6_15 ? 4'hf : _T_89096; // @[LoadQueue.scala 191:60:@38316.4]
  assign _T_89100 = conflictPReg_6_0 | conflictPReg_6_1; // @[LoadQueue.scala 192:43:@38318.4]
  assign _T_89101 = _T_89100 | conflictPReg_6_2; // @[LoadQueue.scala 192:43:@38319.4]
  assign _T_89102 = _T_89101 | conflictPReg_6_3; // @[LoadQueue.scala 192:43:@38320.4]
  assign _T_89103 = _T_89102 | conflictPReg_6_4; // @[LoadQueue.scala 192:43:@38321.4]
  assign _T_89104 = _T_89103 | conflictPReg_6_5; // @[LoadQueue.scala 192:43:@38322.4]
  assign _T_89105 = _T_89104 | conflictPReg_6_6; // @[LoadQueue.scala 192:43:@38323.4]
  assign _T_89106 = _T_89105 | conflictPReg_6_7; // @[LoadQueue.scala 192:43:@38324.4]
  assign _T_89107 = _T_89106 | conflictPReg_6_8; // @[LoadQueue.scala 192:43:@38325.4]
  assign _T_89108 = _T_89107 | conflictPReg_6_9; // @[LoadQueue.scala 192:43:@38326.4]
  assign _T_89109 = _T_89108 | conflictPReg_6_10; // @[LoadQueue.scala 192:43:@38327.4]
  assign _T_89110 = _T_89109 | conflictPReg_6_11; // @[LoadQueue.scala 192:43:@38328.4]
  assign _T_89111 = _T_89110 | conflictPReg_6_12; // @[LoadQueue.scala 192:43:@38329.4]
  assign _T_89112 = _T_89111 | conflictPReg_6_13; // @[LoadQueue.scala 192:43:@38330.4]
  assign _T_89113 = _T_89112 | conflictPReg_6_14; // @[LoadQueue.scala 192:43:@38331.4]
  assign _T_89114 = _T_89113 | conflictPReg_6_15; // @[LoadQueue.scala 192:43:@38332.4]
  assign _GEN_1260 = 4'h0 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1261 = 4'h1 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1262 = 4'h2 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1263 = 4'h3 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1264 = 4'h4 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1265 = 4'h5 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1266 = 4'h6 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1267 = 4'h7 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1268 = 4'h8 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1269 = 4'h9 == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1270 = 4'ha == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1271 = 4'hb == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1272 = 4'hc == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1273 = 4'hd == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1274 = 4'he == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1275 = 4'hf == _T_89097; // @[LoadQueue.scala 193:43:@38334.6]
  assign _GEN_1277 = 4'h1 == _T_89097 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1278 = 4'h2 == _T_89097 ? shiftedStoreDataKnownPReg_2 : _GEN_1277; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1279 = 4'h3 == _T_89097 ? shiftedStoreDataKnownPReg_3 : _GEN_1278; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1280 = 4'h4 == _T_89097 ? shiftedStoreDataKnownPReg_4 : _GEN_1279; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1281 = 4'h5 == _T_89097 ? shiftedStoreDataKnownPReg_5 : _GEN_1280; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1282 = 4'h6 == _T_89097 ? shiftedStoreDataKnownPReg_6 : _GEN_1281; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1283 = 4'h7 == _T_89097 ? shiftedStoreDataKnownPReg_7 : _GEN_1282; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1284 = 4'h8 == _T_89097 ? shiftedStoreDataKnownPReg_8 : _GEN_1283; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1285 = 4'h9 == _T_89097 ? shiftedStoreDataKnownPReg_9 : _GEN_1284; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1286 = 4'ha == _T_89097 ? shiftedStoreDataKnownPReg_10 : _GEN_1285; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1287 = 4'hb == _T_89097 ? shiftedStoreDataKnownPReg_11 : _GEN_1286; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1288 = 4'hc == _T_89097 ? shiftedStoreDataKnownPReg_12 : _GEN_1287; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1289 = 4'hd == _T_89097 ? shiftedStoreDataKnownPReg_13 : _GEN_1288; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1290 = 4'he == _T_89097 ? shiftedStoreDataKnownPReg_14 : _GEN_1289; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1291 = 4'hf == _T_89097 ? shiftedStoreDataKnownPReg_15 : _GEN_1290; // @[LoadQueue.scala 194:31:@38335.6]
  assign _GEN_1293 = 4'h1 == _T_89097 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1294 = 4'h2 == _T_89097 ? shiftedStoreDataQPreg_2 : _GEN_1293; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1295 = 4'h3 == _T_89097 ? shiftedStoreDataQPreg_3 : _GEN_1294; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1296 = 4'h4 == _T_89097 ? shiftedStoreDataQPreg_4 : _GEN_1295; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1297 = 4'h5 == _T_89097 ? shiftedStoreDataQPreg_5 : _GEN_1296; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1298 = 4'h6 == _T_89097 ? shiftedStoreDataQPreg_6 : _GEN_1297; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1299 = 4'h7 == _T_89097 ? shiftedStoreDataQPreg_7 : _GEN_1298; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1300 = 4'h8 == _T_89097 ? shiftedStoreDataQPreg_8 : _GEN_1299; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1301 = 4'h9 == _T_89097 ? shiftedStoreDataQPreg_9 : _GEN_1300; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1302 = 4'ha == _T_89097 ? shiftedStoreDataQPreg_10 : _GEN_1301; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1303 = 4'hb == _T_89097 ? shiftedStoreDataQPreg_11 : _GEN_1302; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1304 = 4'hc == _T_89097 ? shiftedStoreDataQPreg_12 : _GEN_1303; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1305 = 4'hd == _T_89097 ? shiftedStoreDataQPreg_13 : _GEN_1304; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1306 = 4'he == _T_89097 ? shiftedStoreDataQPreg_14 : _GEN_1305; // @[LoadQueue.scala 195:31:@38336.6]
  assign _GEN_1307 = 4'hf == _T_89097 ? shiftedStoreDataQPreg_15 : _GEN_1306; // @[LoadQueue.scala 195:31:@38336.6]
  assign lastConflict_6_0 = _T_89114 ? _GEN_1260 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_1 = _T_89114 ? _GEN_1261 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_2 = _T_89114 ? _GEN_1262 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_3 = _T_89114 ? _GEN_1263 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_4 = _T_89114 ? _GEN_1264 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_5 = _T_89114 ? _GEN_1265 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_6 = _T_89114 ? _GEN_1266 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_7 = _T_89114 ? _GEN_1267 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_8 = _T_89114 ? _GEN_1268 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_9 = _T_89114 ? _GEN_1269 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_10 = _T_89114 ? _GEN_1270 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_11 = _T_89114 ? _GEN_1271 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_12 = _T_89114 ? _GEN_1272 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_13 = _T_89114 ? _GEN_1273 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_14 = _T_89114 ? _GEN_1274 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign lastConflict_6_15 = _T_89114 ? _GEN_1275 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign canBypass_6 = _T_89114 ? _GEN_1291 : 1'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign bypassVal_6 = _T_89114 ? _GEN_1307 : 32'h0; // @[LoadQueue.scala 192:53:@38333.4]
  assign _T_89220 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[LoadQueue.scala 191:60:@38390.4]
  assign _T_89221 = conflictPReg_7_3 ? 2'h3 : _T_89220; // @[LoadQueue.scala 191:60:@38391.4]
  assign _T_89222 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_89221}; // @[LoadQueue.scala 191:60:@38392.4]
  assign _T_89223 = conflictPReg_7_5 ? 3'h5 : _T_89222; // @[LoadQueue.scala 191:60:@38393.4]
  assign _T_89224 = conflictPReg_7_6 ? 3'h6 : _T_89223; // @[LoadQueue.scala 191:60:@38394.4]
  assign _T_89225 = conflictPReg_7_7 ? 3'h7 : _T_89224; // @[LoadQueue.scala 191:60:@38395.4]
  assign _T_89226 = conflictPReg_7_8 ? 4'h8 : {{1'd0}, _T_89225}; // @[LoadQueue.scala 191:60:@38396.4]
  assign _T_89227 = conflictPReg_7_9 ? 4'h9 : _T_89226; // @[LoadQueue.scala 191:60:@38397.4]
  assign _T_89228 = conflictPReg_7_10 ? 4'ha : _T_89227; // @[LoadQueue.scala 191:60:@38398.4]
  assign _T_89229 = conflictPReg_7_11 ? 4'hb : _T_89228; // @[LoadQueue.scala 191:60:@38399.4]
  assign _T_89230 = conflictPReg_7_12 ? 4'hc : _T_89229; // @[LoadQueue.scala 191:60:@38400.4]
  assign _T_89231 = conflictPReg_7_13 ? 4'hd : _T_89230; // @[LoadQueue.scala 191:60:@38401.4]
  assign _T_89232 = conflictPReg_7_14 ? 4'he : _T_89231; // @[LoadQueue.scala 191:60:@38402.4]
  assign _T_89233 = conflictPReg_7_15 ? 4'hf : _T_89232; // @[LoadQueue.scala 191:60:@38403.4]
  assign _T_89236 = conflictPReg_7_0 | conflictPReg_7_1; // @[LoadQueue.scala 192:43:@38405.4]
  assign _T_89237 = _T_89236 | conflictPReg_7_2; // @[LoadQueue.scala 192:43:@38406.4]
  assign _T_89238 = _T_89237 | conflictPReg_7_3; // @[LoadQueue.scala 192:43:@38407.4]
  assign _T_89239 = _T_89238 | conflictPReg_7_4; // @[LoadQueue.scala 192:43:@38408.4]
  assign _T_89240 = _T_89239 | conflictPReg_7_5; // @[LoadQueue.scala 192:43:@38409.4]
  assign _T_89241 = _T_89240 | conflictPReg_7_6; // @[LoadQueue.scala 192:43:@38410.4]
  assign _T_89242 = _T_89241 | conflictPReg_7_7; // @[LoadQueue.scala 192:43:@38411.4]
  assign _T_89243 = _T_89242 | conflictPReg_7_8; // @[LoadQueue.scala 192:43:@38412.4]
  assign _T_89244 = _T_89243 | conflictPReg_7_9; // @[LoadQueue.scala 192:43:@38413.4]
  assign _T_89245 = _T_89244 | conflictPReg_7_10; // @[LoadQueue.scala 192:43:@38414.4]
  assign _T_89246 = _T_89245 | conflictPReg_7_11; // @[LoadQueue.scala 192:43:@38415.4]
  assign _T_89247 = _T_89246 | conflictPReg_7_12; // @[LoadQueue.scala 192:43:@38416.4]
  assign _T_89248 = _T_89247 | conflictPReg_7_13; // @[LoadQueue.scala 192:43:@38417.4]
  assign _T_89249 = _T_89248 | conflictPReg_7_14; // @[LoadQueue.scala 192:43:@38418.4]
  assign _T_89250 = _T_89249 | conflictPReg_7_15; // @[LoadQueue.scala 192:43:@38419.4]
  assign _GEN_1326 = 4'h0 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1327 = 4'h1 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1328 = 4'h2 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1329 = 4'h3 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1330 = 4'h4 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1331 = 4'h5 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1332 = 4'h6 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1333 = 4'h7 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1334 = 4'h8 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1335 = 4'h9 == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1336 = 4'ha == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1337 = 4'hb == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1338 = 4'hc == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1339 = 4'hd == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1340 = 4'he == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1341 = 4'hf == _T_89233; // @[LoadQueue.scala 193:43:@38421.6]
  assign _GEN_1343 = 4'h1 == _T_89233 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1344 = 4'h2 == _T_89233 ? shiftedStoreDataKnownPReg_2 : _GEN_1343; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1345 = 4'h3 == _T_89233 ? shiftedStoreDataKnownPReg_3 : _GEN_1344; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1346 = 4'h4 == _T_89233 ? shiftedStoreDataKnownPReg_4 : _GEN_1345; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1347 = 4'h5 == _T_89233 ? shiftedStoreDataKnownPReg_5 : _GEN_1346; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1348 = 4'h6 == _T_89233 ? shiftedStoreDataKnownPReg_6 : _GEN_1347; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1349 = 4'h7 == _T_89233 ? shiftedStoreDataKnownPReg_7 : _GEN_1348; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1350 = 4'h8 == _T_89233 ? shiftedStoreDataKnownPReg_8 : _GEN_1349; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1351 = 4'h9 == _T_89233 ? shiftedStoreDataKnownPReg_9 : _GEN_1350; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1352 = 4'ha == _T_89233 ? shiftedStoreDataKnownPReg_10 : _GEN_1351; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1353 = 4'hb == _T_89233 ? shiftedStoreDataKnownPReg_11 : _GEN_1352; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1354 = 4'hc == _T_89233 ? shiftedStoreDataKnownPReg_12 : _GEN_1353; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1355 = 4'hd == _T_89233 ? shiftedStoreDataKnownPReg_13 : _GEN_1354; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1356 = 4'he == _T_89233 ? shiftedStoreDataKnownPReg_14 : _GEN_1355; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1357 = 4'hf == _T_89233 ? shiftedStoreDataKnownPReg_15 : _GEN_1356; // @[LoadQueue.scala 194:31:@38422.6]
  assign _GEN_1359 = 4'h1 == _T_89233 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1360 = 4'h2 == _T_89233 ? shiftedStoreDataQPreg_2 : _GEN_1359; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1361 = 4'h3 == _T_89233 ? shiftedStoreDataQPreg_3 : _GEN_1360; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1362 = 4'h4 == _T_89233 ? shiftedStoreDataQPreg_4 : _GEN_1361; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1363 = 4'h5 == _T_89233 ? shiftedStoreDataQPreg_5 : _GEN_1362; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1364 = 4'h6 == _T_89233 ? shiftedStoreDataQPreg_6 : _GEN_1363; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1365 = 4'h7 == _T_89233 ? shiftedStoreDataQPreg_7 : _GEN_1364; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1366 = 4'h8 == _T_89233 ? shiftedStoreDataQPreg_8 : _GEN_1365; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1367 = 4'h9 == _T_89233 ? shiftedStoreDataQPreg_9 : _GEN_1366; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1368 = 4'ha == _T_89233 ? shiftedStoreDataQPreg_10 : _GEN_1367; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1369 = 4'hb == _T_89233 ? shiftedStoreDataQPreg_11 : _GEN_1368; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1370 = 4'hc == _T_89233 ? shiftedStoreDataQPreg_12 : _GEN_1369; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1371 = 4'hd == _T_89233 ? shiftedStoreDataQPreg_13 : _GEN_1370; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1372 = 4'he == _T_89233 ? shiftedStoreDataQPreg_14 : _GEN_1371; // @[LoadQueue.scala 195:31:@38423.6]
  assign _GEN_1373 = 4'hf == _T_89233 ? shiftedStoreDataQPreg_15 : _GEN_1372; // @[LoadQueue.scala 195:31:@38423.6]
  assign lastConflict_7_0 = _T_89250 ? _GEN_1326 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_1 = _T_89250 ? _GEN_1327 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_2 = _T_89250 ? _GEN_1328 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_3 = _T_89250 ? _GEN_1329 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_4 = _T_89250 ? _GEN_1330 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_5 = _T_89250 ? _GEN_1331 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_6 = _T_89250 ? _GEN_1332 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_7 = _T_89250 ? _GEN_1333 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_8 = _T_89250 ? _GEN_1334 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_9 = _T_89250 ? _GEN_1335 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_10 = _T_89250 ? _GEN_1336 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_11 = _T_89250 ? _GEN_1337 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_12 = _T_89250 ? _GEN_1338 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_13 = _T_89250 ? _GEN_1339 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_14 = _T_89250 ? _GEN_1340 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign lastConflict_7_15 = _T_89250 ? _GEN_1341 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign canBypass_7 = _T_89250 ? _GEN_1357 : 1'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign bypassVal_7 = _T_89250 ? _GEN_1373 : 32'h0; // @[LoadQueue.scala 192:53:@38420.4]
  assign _T_89356 = conflictPReg_8_2 ? 2'h2 : {{1'd0}, conflictPReg_8_1}; // @[LoadQueue.scala 191:60:@38477.4]
  assign _T_89357 = conflictPReg_8_3 ? 2'h3 : _T_89356; // @[LoadQueue.scala 191:60:@38478.4]
  assign _T_89358 = conflictPReg_8_4 ? 3'h4 : {{1'd0}, _T_89357}; // @[LoadQueue.scala 191:60:@38479.4]
  assign _T_89359 = conflictPReg_8_5 ? 3'h5 : _T_89358; // @[LoadQueue.scala 191:60:@38480.4]
  assign _T_89360 = conflictPReg_8_6 ? 3'h6 : _T_89359; // @[LoadQueue.scala 191:60:@38481.4]
  assign _T_89361 = conflictPReg_8_7 ? 3'h7 : _T_89360; // @[LoadQueue.scala 191:60:@38482.4]
  assign _T_89362 = conflictPReg_8_8 ? 4'h8 : {{1'd0}, _T_89361}; // @[LoadQueue.scala 191:60:@38483.4]
  assign _T_89363 = conflictPReg_8_9 ? 4'h9 : _T_89362; // @[LoadQueue.scala 191:60:@38484.4]
  assign _T_89364 = conflictPReg_8_10 ? 4'ha : _T_89363; // @[LoadQueue.scala 191:60:@38485.4]
  assign _T_89365 = conflictPReg_8_11 ? 4'hb : _T_89364; // @[LoadQueue.scala 191:60:@38486.4]
  assign _T_89366 = conflictPReg_8_12 ? 4'hc : _T_89365; // @[LoadQueue.scala 191:60:@38487.4]
  assign _T_89367 = conflictPReg_8_13 ? 4'hd : _T_89366; // @[LoadQueue.scala 191:60:@38488.4]
  assign _T_89368 = conflictPReg_8_14 ? 4'he : _T_89367; // @[LoadQueue.scala 191:60:@38489.4]
  assign _T_89369 = conflictPReg_8_15 ? 4'hf : _T_89368; // @[LoadQueue.scala 191:60:@38490.4]
  assign _T_89372 = conflictPReg_8_0 | conflictPReg_8_1; // @[LoadQueue.scala 192:43:@38492.4]
  assign _T_89373 = _T_89372 | conflictPReg_8_2; // @[LoadQueue.scala 192:43:@38493.4]
  assign _T_89374 = _T_89373 | conflictPReg_8_3; // @[LoadQueue.scala 192:43:@38494.4]
  assign _T_89375 = _T_89374 | conflictPReg_8_4; // @[LoadQueue.scala 192:43:@38495.4]
  assign _T_89376 = _T_89375 | conflictPReg_8_5; // @[LoadQueue.scala 192:43:@38496.4]
  assign _T_89377 = _T_89376 | conflictPReg_8_6; // @[LoadQueue.scala 192:43:@38497.4]
  assign _T_89378 = _T_89377 | conflictPReg_8_7; // @[LoadQueue.scala 192:43:@38498.4]
  assign _T_89379 = _T_89378 | conflictPReg_8_8; // @[LoadQueue.scala 192:43:@38499.4]
  assign _T_89380 = _T_89379 | conflictPReg_8_9; // @[LoadQueue.scala 192:43:@38500.4]
  assign _T_89381 = _T_89380 | conflictPReg_8_10; // @[LoadQueue.scala 192:43:@38501.4]
  assign _T_89382 = _T_89381 | conflictPReg_8_11; // @[LoadQueue.scala 192:43:@38502.4]
  assign _T_89383 = _T_89382 | conflictPReg_8_12; // @[LoadQueue.scala 192:43:@38503.4]
  assign _T_89384 = _T_89383 | conflictPReg_8_13; // @[LoadQueue.scala 192:43:@38504.4]
  assign _T_89385 = _T_89384 | conflictPReg_8_14; // @[LoadQueue.scala 192:43:@38505.4]
  assign _T_89386 = _T_89385 | conflictPReg_8_15; // @[LoadQueue.scala 192:43:@38506.4]
  assign _GEN_1392 = 4'h0 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1393 = 4'h1 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1394 = 4'h2 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1395 = 4'h3 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1396 = 4'h4 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1397 = 4'h5 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1398 = 4'h6 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1399 = 4'h7 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1400 = 4'h8 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1401 = 4'h9 == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1402 = 4'ha == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1403 = 4'hb == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1404 = 4'hc == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1405 = 4'hd == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1406 = 4'he == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1407 = 4'hf == _T_89369; // @[LoadQueue.scala 193:43:@38508.6]
  assign _GEN_1409 = 4'h1 == _T_89369 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1410 = 4'h2 == _T_89369 ? shiftedStoreDataKnownPReg_2 : _GEN_1409; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1411 = 4'h3 == _T_89369 ? shiftedStoreDataKnownPReg_3 : _GEN_1410; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1412 = 4'h4 == _T_89369 ? shiftedStoreDataKnownPReg_4 : _GEN_1411; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1413 = 4'h5 == _T_89369 ? shiftedStoreDataKnownPReg_5 : _GEN_1412; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1414 = 4'h6 == _T_89369 ? shiftedStoreDataKnownPReg_6 : _GEN_1413; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1415 = 4'h7 == _T_89369 ? shiftedStoreDataKnownPReg_7 : _GEN_1414; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1416 = 4'h8 == _T_89369 ? shiftedStoreDataKnownPReg_8 : _GEN_1415; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1417 = 4'h9 == _T_89369 ? shiftedStoreDataKnownPReg_9 : _GEN_1416; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1418 = 4'ha == _T_89369 ? shiftedStoreDataKnownPReg_10 : _GEN_1417; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1419 = 4'hb == _T_89369 ? shiftedStoreDataKnownPReg_11 : _GEN_1418; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1420 = 4'hc == _T_89369 ? shiftedStoreDataKnownPReg_12 : _GEN_1419; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1421 = 4'hd == _T_89369 ? shiftedStoreDataKnownPReg_13 : _GEN_1420; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1422 = 4'he == _T_89369 ? shiftedStoreDataKnownPReg_14 : _GEN_1421; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1423 = 4'hf == _T_89369 ? shiftedStoreDataKnownPReg_15 : _GEN_1422; // @[LoadQueue.scala 194:31:@38509.6]
  assign _GEN_1425 = 4'h1 == _T_89369 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1426 = 4'h2 == _T_89369 ? shiftedStoreDataQPreg_2 : _GEN_1425; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1427 = 4'h3 == _T_89369 ? shiftedStoreDataQPreg_3 : _GEN_1426; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1428 = 4'h4 == _T_89369 ? shiftedStoreDataQPreg_4 : _GEN_1427; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1429 = 4'h5 == _T_89369 ? shiftedStoreDataQPreg_5 : _GEN_1428; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1430 = 4'h6 == _T_89369 ? shiftedStoreDataQPreg_6 : _GEN_1429; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1431 = 4'h7 == _T_89369 ? shiftedStoreDataQPreg_7 : _GEN_1430; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1432 = 4'h8 == _T_89369 ? shiftedStoreDataQPreg_8 : _GEN_1431; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1433 = 4'h9 == _T_89369 ? shiftedStoreDataQPreg_9 : _GEN_1432; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1434 = 4'ha == _T_89369 ? shiftedStoreDataQPreg_10 : _GEN_1433; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1435 = 4'hb == _T_89369 ? shiftedStoreDataQPreg_11 : _GEN_1434; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1436 = 4'hc == _T_89369 ? shiftedStoreDataQPreg_12 : _GEN_1435; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1437 = 4'hd == _T_89369 ? shiftedStoreDataQPreg_13 : _GEN_1436; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1438 = 4'he == _T_89369 ? shiftedStoreDataQPreg_14 : _GEN_1437; // @[LoadQueue.scala 195:31:@38510.6]
  assign _GEN_1439 = 4'hf == _T_89369 ? shiftedStoreDataQPreg_15 : _GEN_1438; // @[LoadQueue.scala 195:31:@38510.6]
  assign lastConflict_8_0 = _T_89386 ? _GEN_1392 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_1 = _T_89386 ? _GEN_1393 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_2 = _T_89386 ? _GEN_1394 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_3 = _T_89386 ? _GEN_1395 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_4 = _T_89386 ? _GEN_1396 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_5 = _T_89386 ? _GEN_1397 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_6 = _T_89386 ? _GEN_1398 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_7 = _T_89386 ? _GEN_1399 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_8 = _T_89386 ? _GEN_1400 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_9 = _T_89386 ? _GEN_1401 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_10 = _T_89386 ? _GEN_1402 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_11 = _T_89386 ? _GEN_1403 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_12 = _T_89386 ? _GEN_1404 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_13 = _T_89386 ? _GEN_1405 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_14 = _T_89386 ? _GEN_1406 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign lastConflict_8_15 = _T_89386 ? _GEN_1407 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign canBypass_8 = _T_89386 ? _GEN_1423 : 1'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign bypassVal_8 = _T_89386 ? _GEN_1439 : 32'h0; // @[LoadQueue.scala 192:53:@38507.4]
  assign _T_89492 = conflictPReg_9_2 ? 2'h2 : {{1'd0}, conflictPReg_9_1}; // @[LoadQueue.scala 191:60:@38564.4]
  assign _T_89493 = conflictPReg_9_3 ? 2'h3 : _T_89492; // @[LoadQueue.scala 191:60:@38565.4]
  assign _T_89494 = conflictPReg_9_4 ? 3'h4 : {{1'd0}, _T_89493}; // @[LoadQueue.scala 191:60:@38566.4]
  assign _T_89495 = conflictPReg_9_5 ? 3'h5 : _T_89494; // @[LoadQueue.scala 191:60:@38567.4]
  assign _T_89496 = conflictPReg_9_6 ? 3'h6 : _T_89495; // @[LoadQueue.scala 191:60:@38568.4]
  assign _T_89497 = conflictPReg_9_7 ? 3'h7 : _T_89496; // @[LoadQueue.scala 191:60:@38569.4]
  assign _T_89498 = conflictPReg_9_8 ? 4'h8 : {{1'd0}, _T_89497}; // @[LoadQueue.scala 191:60:@38570.4]
  assign _T_89499 = conflictPReg_9_9 ? 4'h9 : _T_89498; // @[LoadQueue.scala 191:60:@38571.4]
  assign _T_89500 = conflictPReg_9_10 ? 4'ha : _T_89499; // @[LoadQueue.scala 191:60:@38572.4]
  assign _T_89501 = conflictPReg_9_11 ? 4'hb : _T_89500; // @[LoadQueue.scala 191:60:@38573.4]
  assign _T_89502 = conflictPReg_9_12 ? 4'hc : _T_89501; // @[LoadQueue.scala 191:60:@38574.4]
  assign _T_89503 = conflictPReg_9_13 ? 4'hd : _T_89502; // @[LoadQueue.scala 191:60:@38575.4]
  assign _T_89504 = conflictPReg_9_14 ? 4'he : _T_89503; // @[LoadQueue.scala 191:60:@38576.4]
  assign _T_89505 = conflictPReg_9_15 ? 4'hf : _T_89504; // @[LoadQueue.scala 191:60:@38577.4]
  assign _T_89508 = conflictPReg_9_0 | conflictPReg_9_1; // @[LoadQueue.scala 192:43:@38579.4]
  assign _T_89509 = _T_89508 | conflictPReg_9_2; // @[LoadQueue.scala 192:43:@38580.4]
  assign _T_89510 = _T_89509 | conflictPReg_9_3; // @[LoadQueue.scala 192:43:@38581.4]
  assign _T_89511 = _T_89510 | conflictPReg_9_4; // @[LoadQueue.scala 192:43:@38582.4]
  assign _T_89512 = _T_89511 | conflictPReg_9_5; // @[LoadQueue.scala 192:43:@38583.4]
  assign _T_89513 = _T_89512 | conflictPReg_9_6; // @[LoadQueue.scala 192:43:@38584.4]
  assign _T_89514 = _T_89513 | conflictPReg_9_7; // @[LoadQueue.scala 192:43:@38585.4]
  assign _T_89515 = _T_89514 | conflictPReg_9_8; // @[LoadQueue.scala 192:43:@38586.4]
  assign _T_89516 = _T_89515 | conflictPReg_9_9; // @[LoadQueue.scala 192:43:@38587.4]
  assign _T_89517 = _T_89516 | conflictPReg_9_10; // @[LoadQueue.scala 192:43:@38588.4]
  assign _T_89518 = _T_89517 | conflictPReg_9_11; // @[LoadQueue.scala 192:43:@38589.4]
  assign _T_89519 = _T_89518 | conflictPReg_9_12; // @[LoadQueue.scala 192:43:@38590.4]
  assign _T_89520 = _T_89519 | conflictPReg_9_13; // @[LoadQueue.scala 192:43:@38591.4]
  assign _T_89521 = _T_89520 | conflictPReg_9_14; // @[LoadQueue.scala 192:43:@38592.4]
  assign _T_89522 = _T_89521 | conflictPReg_9_15; // @[LoadQueue.scala 192:43:@38593.4]
  assign _GEN_1458 = 4'h0 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1459 = 4'h1 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1460 = 4'h2 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1461 = 4'h3 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1462 = 4'h4 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1463 = 4'h5 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1464 = 4'h6 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1465 = 4'h7 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1466 = 4'h8 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1467 = 4'h9 == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1468 = 4'ha == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1469 = 4'hb == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1470 = 4'hc == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1471 = 4'hd == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1472 = 4'he == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1473 = 4'hf == _T_89505; // @[LoadQueue.scala 193:43:@38595.6]
  assign _GEN_1475 = 4'h1 == _T_89505 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1476 = 4'h2 == _T_89505 ? shiftedStoreDataKnownPReg_2 : _GEN_1475; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1477 = 4'h3 == _T_89505 ? shiftedStoreDataKnownPReg_3 : _GEN_1476; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1478 = 4'h4 == _T_89505 ? shiftedStoreDataKnownPReg_4 : _GEN_1477; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1479 = 4'h5 == _T_89505 ? shiftedStoreDataKnownPReg_5 : _GEN_1478; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1480 = 4'h6 == _T_89505 ? shiftedStoreDataKnownPReg_6 : _GEN_1479; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1481 = 4'h7 == _T_89505 ? shiftedStoreDataKnownPReg_7 : _GEN_1480; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1482 = 4'h8 == _T_89505 ? shiftedStoreDataKnownPReg_8 : _GEN_1481; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1483 = 4'h9 == _T_89505 ? shiftedStoreDataKnownPReg_9 : _GEN_1482; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1484 = 4'ha == _T_89505 ? shiftedStoreDataKnownPReg_10 : _GEN_1483; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1485 = 4'hb == _T_89505 ? shiftedStoreDataKnownPReg_11 : _GEN_1484; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1486 = 4'hc == _T_89505 ? shiftedStoreDataKnownPReg_12 : _GEN_1485; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1487 = 4'hd == _T_89505 ? shiftedStoreDataKnownPReg_13 : _GEN_1486; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1488 = 4'he == _T_89505 ? shiftedStoreDataKnownPReg_14 : _GEN_1487; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1489 = 4'hf == _T_89505 ? shiftedStoreDataKnownPReg_15 : _GEN_1488; // @[LoadQueue.scala 194:31:@38596.6]
  assign _GEN_1491 = 4'h1 == _T_89505 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1492 = 4'h2 == _T_89505 ? shiftedStoreDataQPreg_2 : _GEN_1491; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1493 = 4'h3 == _T_89505 ? shiftedStoreDataQPreg_3 : _GEN_1492; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1494 = 4'h4 == _T_89505 ? shiftedStoreDataQPreg_4 : _GEN_1493; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1495 = 4'h5 == _T_89505 ? shiftedStoreDataQPreg_5 : _GEN_1494; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1496 = 4'h6 == _T_89505 ? shiftedStoreDataQPreg_6 : _GEN_1495; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1497 = 4'h7 == _T_89505 ? shiftedStoreDataQPreg_7 : _GEN_1496; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1498 = 4'h8 == _T_89505 ? shiftedStoreDataQPreg_8 : _GEN_1497; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1499 = 4'h9 == _T_89505 ? shiftedStoreDataQPreg_9 : _GEN_1498; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1500 = 4'ha == _T_89505 ? shiftedStoreDataQPreg_10 : _GEN_1499; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1501 = 4'hb == _T_89505 ? shiftedStoreDataQPreg_11 : _GEN_1500; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1502 = 4'hc == _T_89505 ? shiftedStoreDataQPreg_12 : _GEN_1501; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1503 = 4'hd == _T_89505 ? shiftedStoreDataQPreg_13 : _GEN_1502; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1504 = 4'he == _T_89505 ? shiftedStoreDataQPreg_14 : _GEN_1503; // @[LoadQueue.scala 195:31:@38597.6]
  assign _GEN_1505 = 4'hf == _T_89505 ? shiftedStoreDataQPreg_15 : _GEN_1504; // @[LoadQueue.scala 195:31:@38597.6]
  assign lastConflict_9_0 = _T_89522 ? _GEN_1458 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_1 = _T_89522 ? _GEN_1459 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_2 = _T_89522 ? _GEN_1460 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_3 = _T_89522 ? _GEN_1461 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_4 = _T_89522 ? _GEN_1462 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_5 = _T_89522 ? _GEN_1463 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_6 = _T_89522 ? _GEN_1464 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_7 = _T_89522 ? _GEN_1465 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_8 = _T_89522 ? _GEN_1466 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_9 = _T_89522 ? _GEN_1467 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_10 = _T_89522 ? _GEN_1468 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_11 = _T_89522 ? _GEN_1469 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_12 = _T_89522 ? _GEN_1470 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_13 = _T_89522 ? _GEN_1471 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_14 = _T_89522 ? _GEN_1472 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign lastConflict_9_15 = _T_89522 ? _GEN_1473 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign canBypass_9 = _T_89522 ? _GEN_1489 : 1'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign bypassVal_9 = _T_89522 ? _GEN_1505 : 32'h0; // @[LoadQueue.scala 192:53:@38594.4]
  assign _T_89628 = conflictPReg_10_2 ? 2'h2 : {{1'd0}, conflictPReg_10_1}; // @[LoadQueue.scala 191:60:@38651.4]
  assign _T_89629 = conflictPReg_10_3 ? 2'h3 : _T_89628; // @[LoadQueue.scala 191:60:@38652.4]
  assign _T_89630 = conflictPReg_10_4 ? 3'h4 : {{1'd0}, _T_89629}; // @[LoadQueue.scala 191:60:@38653.4]
  assign _T_89631 = conflictPReg_10_5 ? 3'h5 : _T_89630; // @[LoadQueue.scala 191:60:@38654.4]
  assign _T_89632 = conflictPReg_10_6 ? 3'h6 : _T_89631; // @[LoadQueue.scala 191:60:@38655.4]
  assign _T_89633 = conflictPReg_10_7 ? 3'h7 : _T_89632; // @[LoadQueue.scala 191:60:@38656.4]
  assign _T_89634 = conflictPReg_10_8 ? 4'h8 : {{1'd0}, _T_89633}; // @[LoadQueue.scala 191:60:@38657.4]
  assign _T_89635 = conflictPReg_10_9 ? 4'h9 : _T_89634; // @[LoadQueue.scala 191:60:@38658.4]
  assign _T_89636 = conflictPReg_10_10 ? 4'ha : _T_89635; // @[LoadQueue.scala 191:60:@38659.4]
  assign _T_89637 = conflictPReg_10_11 ? 4'hb : _T_89636; // @[LoadQueue.scala 191:60:@38660.4]
  assign _T_89638 = conflictPReg_10_12 ? 4'hc : _T_89637; // @[LoadQueue.scala 191:60:@38661.4]
  assign _T_89639 = conflictPReg_10_13 ? 4'hd : _T_89638; // @[LoadQueue.scala 191:60:@38662.4]
  assign _T_89640 = conflictPReg_10_14 ? 4'he : _T_89639; // @[LoadQueue.scala 191:60:@38663.4]
  assign _T_89641 = conflictPReg_10_15 ? 4'hf : _T_89640; // @[LoadQueue.scala 191:60:@38664.4]
  assign _T_89644 = conflictPReg_10_0 | conflictPReg_10_1; // @[LoadQueue.scala 192:43:@38666.4]
  assign _T_89645 = _T_89644 | conflictPReg_10_2; // @[LoadQueue.scala 192:43:@38667.4]
  assign _T_89646 = _T_89645 | conflictPReg_10_3; // @[LoadQueue.scala 192:43:@38668.4]
  assign _T_89647 = _T_89646 | conflictPReg_10_4; // @[LoadQueue.scala 192:43:@38669.4]
  assign _T_89648 = _T_89647 | conflictPReg_10_5; // @[LoadQueue.scala 192:43:@38670.4]
  assign _T_89649 = _T_89648 | conflictPReg_10_6; // @[LoadQueue.scala 192:43:@38671.4]
  assign _T_89650 = _T_89649 | conflictPReg_10_7; // @[LoadQueue.scala 192:43:@38672.4]
  assign _T_89651 = _T_89650 | conflictPReg_10_8; // @[LoadQueue.scala 192:43:@38673.4]
  assign _T_89652 = _T_89651 | conflictPReg_10_9; // @[LoadQueue.scala 192:43:@38674.4]
  assign _T_89653 = _T_89652 | conflictPReg_10_10; // @[LoadQueue.scala 192:43:@38675.4]
  assign _T_89654 = _T_89653 | conflictPReg_10_11; // @[LoadQueue.scala 192:43:@38676.4]
  assign _T_89655 = _T_89654 | conflictPReg_10_12; // @[LoadQueue.scala 192:43:@38677.4]
  assign _T_89656 = _T_89655 | conflictPReg_10_13; // @[LoadQueue.scala 192:43:@38678.4]
  assign _T_89657 = _T_89656 | conflictPReg_10_14; // @[LoadQueue.scala 192:43:@38679.4]
  assign _T_89658 = _T_89657 | conflictPReg_10_15; // @[LoadQueue.scala 192:43:@38680.4]
  assign _GEN_1524 = 4'h0 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1525 = 4'h1 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1526 = 4'h2 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1527 = 4'h3 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1528 = 4'h4 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1529 = 4'h5 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1530 = 4'h6 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1531 = 4'h7 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1532 = 4'h8 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1533 = 4'h9 == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1534 = 4'ha == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1535 = 4'hb == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1536 = 4'hc == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1537 = 4'hd == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1538 = 4'he == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1539 = 4'hf == _T_89641; // @[LoadQueue.scala 193:43:@38682.6]
  assign _GEN_1541 = 4'h1 == _T_89641 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1542 = 4'h2 == _T_89641 ? shiftedStoreDataKnownPReg_2 : _GEN_1541; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1543 = 4'h3 == _T_89641 ? shiftedStoreDataKnownPReg_3 : _GEN_1542; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1544 = 4'h4 == _T_89641 ? shiftedStoreDataKnownPReg_4 : _GEN_1543; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1545 = 4'h5 == _T_89641 ? shiftedStoreDataKnownPReg_5 : _GEN_1544; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1546 = 4'h6 == _T_89641 ? shiftedStoreDataKnownPReg_6 : _GEN_1545; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1547 = 4'h7 == _T_89641 ? shiftedStoreDataKnownPReg_7 : _GEN_1546; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1548 = 4'h8 == _T_89641 ? shiftedStoreDataKnownPReg_8 : _GEN_1547; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1549 = 4'h9 == _T_89641 ? shiftedStoreDataKnownPReg_9 : _GEN_1548; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1550 = 4'ha == _T_89641 ? shiftedStoreDataKnownPReg_10 : _GEN_1549; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1551 = 4'hb == _T_89641 ? shiftedStoreDataKnownPReg_11 : _GEN_1550; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1552 = 4'hc == _T_89641 ? shiftedStoreDataKnownPReg_12 : _GEN_1551; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1553 = 4'hd == _T_89641 ? shiftedStoreDataKnownPReg_13 : _GEN_1552; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1554 = 4'he == _T_89641 ? shiftedStoreDataKnownPReg_14 : _GEN_1553; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1555 = 4'hf == _T_89641 ? shiftedStoreDataKnownPReg_15 : _GEN_1554; // @[LoadQueue.scala 194:31:@38683.6]
  assign _GEN_1557 = 4'h1 == _T_89641 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1558 = 4'h2 == _T_89641 ? shiftedStoreDataQPreg_2 : _GEN_1557; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1559 = 4'h3 == _T_89641 ? shiftedStoreDataQPreg_3 : _GEN_1558; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1560 = 4'h4 == _T_89641 ? shiftedStoreDataQPreg_4 : _GEN_1559; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1561 = 4'h5 == _T_89641 ? shiftedStoreDataQPreg_5 : _GEN_1560; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1562 = 4'h6 == _T_89641 ? shiftedStoreDataQPreg_6 : _GEN_1561; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1563 = 4'h7 == _T_89641 ? shiftedStoreDataQPreg_7 : _GEN_1562; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1564 = 4'h8 == _T_89641 ? shiftedStoreDataQPreg_8 : _GEN_1563; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1565 = 4'h9 == _T_89641 ? shiftedStoreDataQPreg_9 : _GEN_1564; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1566 = 4'ha == _T_89641 ? shiftedStoreDataQPreg_10 : _GEN_1565; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1567 = 4'hb == _T_89641 ? shiftedStoreDataQPreg_11 : _GEN_1566; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1568 = 4'hc == _T_89641 ? shiftedStoreDataQPreg_12 : _GEN_1567; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1569 = 4'hd == _T_89641 ? shiftedStoreDataQPreg_13 : _GEN_1568; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1570 = 4'he == _T_89641 ? shiftedStoreDataQPreg_14 : _GEN_1569; // @[LoadQueue.scala 195:31:@38684.6]
  assign _GEN_1571 = 4'hf == _T_89641 ? shiftedStoreDataQPreg_15 : _GEN_1570; // @[LoadQueue.scala 195:31:@38684.6]
  assign lastConflict_10_0 = _T_89658 ? _GEN_1524 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_1 = _T_89658 ? _GEN_1525 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_2 = _T_89658 ? _GEN_1526 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_3 = _T_89658 ? _GEN_1527 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_4 = _T_89658 ? _GEN_1528 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_5 = _T_89658 ? _GEN_1529 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_6 = _T_89658 ? _GEN_1530 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_7 = _T_89658 ? _GEN_1531 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_8 = _T_89658 ? _GEN_1532 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_9 = _T_89658 ? _GEN_1533 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_10 = _T_89658 ? _GEN_1534 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_11 = _T_89658 ? _GEN_1535 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_12 = _T_89658 ? _GEN_1536 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_13 = _T_89658 ? _GEN_1537 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_14 = _T_89658 ? _GEN_1538 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign lastConflict_10_15 = _T_89658 ? _GEN_1539 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign canBypass_10 = _T_89658 ? _GEN_1555 : 1'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign bypassVal_10 = _T_89658 ? _GEN_1571 : 32'h0; // @[LoadQueue.scala 192:53:@38681.4]
  assign _T_89764 = conflictPReg_11_2 ? 2'h2 : {{1'd0}, conflictPReg_11_1}; // @[LoadQueue.scala 191:60:@38738.4]
  assign _T_89765 = conflictPReg_11_3 ? 2'h3 : _T_89764; // @[LoadQueue.scala 191:60:@38739.4]
  assign _T_89766 = conflictPReg_11_4 ? 3'h4 : {{1'd0}, _T_89765}; // @[LoadQueue.scala 191:60:@38740.4]
  assign _T_89767 = conflictPReg_11_5 ? 3'h5 : _T_89766; // @[LoadQueue.scala 191:60:@38741.4]
  assign _T_89768 = conflictPReg_11_6 ? 3'h6 : _T_89767; // @[LoadQueue.scala 191:60:@38742.4]
  assign _T_89769 = conflictPReg_11_7 ? 3'h7 : _T_89768; // @[LoadQueue.scala 191:60:@38743.4]
  assign _T_89770 = conflictPReg_11_8 ? 4'h8 : {{1'd0}, _T_89769}; // @[LoadQueue.scala 191:60:@38744.4]
  assign _T_89771 = conflictPReg_11_9 ? 4'h9 : _T_89770; // @[LoadQueue.scala 191:60:@38745.4]
  assign _T_89772 = conflictPReg_11_10 ? 4'ha : _T_89771; // @[LoadQueue.scala 191:60:@38746.4]
  assign _T_89773 = conflictPReg_11_11 ? 4'hb : _T_89772; // @[LoadQueue.scala 191:60:@38747.4]
  assign _T_89774 = conflictPReg_11_12 ? 4'hc : _T_89773; // @[LoadQueue.scala 191:60:@38748.4]
  assign _T_89775 = conflictPReg_11_13 ? 4'hd : _T_89774; // @[LoadQueue.scala 191:60:@38749.4]
  assign _T_89776 = conflictPReg_11_14 ? 4'he : _T_89775; // @[LoadQueue.scala 191:60:@38750.4]
  assign _T_89777 = conflictPReg_11_15 ? 4'hf : _T_89776; // @[LoadQueue.scala 191:60:@38751.4]
  assign _T_89780 = conflictPReg_11_0 | conflictPReg_11_1; // @[LoadQueue.scala 192:43:@38753.4]
  assign _T_89781 = _T_89780 | conflictPReg_11_2; // @[LoadQueue.scala 192:43:@38754.4]
  assign _T_89782 = _T_89781 | conflictPReg_11_3; // @[LoadQueue.scala 192:43:@38755.4]
  assign _T_89783 = _T_89782 | conflictPReg_11_4; // @[LoadQueue.scala 192:43:@38756.4]
  assign _T_89784 = _T_89783 | conflictPReg_11_5; // @[LoadQueue.scala 192:43:@38757.4]
  assign _T_89785 = _T_89784 | conflictPReg_11_6; // @[LoadQueue.scala 192:43:@38758.4]
  assign _T_89786 = _T_89785 | conflictPReg_11_7; // @[LoadQueue.scala 192:43:@38759.4]
  assign _T_89787 = _T_89786 | conflictPReg_11_8; // @[LoadQueue.scala 192:43:@38760.4]
  assign _T_89788 = _T_89787 | conflictPReg_11_9; // @[LoadQueue.scala 192:43:@38761.4]
  assign _T_89789 = _T_89788 | conflictPReg_11_10; // @[LoadQueue.scala 192:43:@38762.4]
  assign _T_89790 = _T_89789 | conflictPReg_11_11; // @[LoadQueue.scala 192:43:@38763.4]
  assign _T_89791 = _T_89790 | conflictPReg_11_12; // @[LoadQueue.scala 192:43:@38764.4]
  assign _T_89792 = _T_89791 | conflictPReg_11_13; // @[LoadQueue.scala 192:43:@38765.4]
  assign _T_89793 = _T_89792 | conflictPReg_11_14; // @[LoadQueue.scala 192:43:@38766.4]
  assign _T_89794 = _T_89793 | conflictPReg_11_15; // @[LoadQueue.scala 192:43:@38767.4]
  assign _GEN_1590 = 4'h0 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1591 = 4'h1 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1592 = 4'h2 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1593 = 4'h3 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1594 = 4'h4 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1595 = 4'h5 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1596 = 4'h6 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1597 = 4'h7 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1598 = 4'h8 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1599 = 4'h9 == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1600 = 4'ha == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1601 = 4'hb == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1602 = 4'hc == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1603 = 4'hd == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1604 = 4'he == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1605 = 4'hf == _T_89777; // @[LoadQueue.scala 193:43:@38769.6]
  assign _GEN_1607 = 4'h1 == _T_89777 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1608 = 4'h2 == _T_89777 ? shiftedStoreDataKnownPReg_2 : _GEN_1607; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1609 = 4'h3 == _T_89777 ? shiftedStoreDataKnownPReg_3 : _GEN_1608; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1610 = 4'h4 == _T_89777 ? shiftedStoreDataKnownPReg_4 : _GEN_1609; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1611 = 4'h5 == _T_89777 ? shiftedStoreDataKnownPReg_5 : _GEN_1610; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1612 = 4'h6 == _T_89777 ? shiftedStoreDataKnownPReg_6 : _GEN_1611; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1613 = 4'h7 == _T_89777 ? shiftedStoreDataKnownPReg_7 : _GEN_1612; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1614 = 4'h8 == _T_89777 ? shiftedStoreDataKnownPReg_8 : _GEN_1613; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1615 = 4'h9 == _T_89777 ? shiftedStoreDataKnownPReg_9 : _GEN_1614; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1616 = 4'ha == _T_89777 ? shiftedStoreDataKnownPReg_10 : _GEN_1615; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1617 = 4'hb == _T_89777 ? shiftedStoreDataKnownPReg_11 : _GEN_1616; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1618 = 4'hc == _T_89777 ? shiftedStoreDataKnownPReg_12 : _GEN_1617; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1619 = 4'hd == _T_89777 ? shiftedStoreDataKnownPReg_13 : _GEN_1618; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1620 = 4'he == _T_89777 ? shiftedStoreDataKnownPReg_14 : _GEN_1619; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1621 = 4'hf == _T_89777 ? shiftedStoreDataKnownPReg_15 : _GEN_1620; // @[LoadQueue.scala 194:31:@38770.6]
  assign _GEN_1623 = 4'h1 == _T_89777 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1624 = 4'h2 == _T_89777 ? shiftedStoreDataQPreg_2 : _GEN_1623; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1625 = 4'h3 == _T_89777 ? shiftedStoreDataQPreg_3 : _GEN_1624; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1626 = 4'h4 == _T_89777 ? shiftedStoreDataQPreg_4 : _GEN_1625; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1627 = 4'h5 == _T_89777 ? shiftedStoreDataQPreg_5 : _GEN_1626; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1628 = 4'h6 == _T_89777 ? shiftedStoreDataQPreg_6 : _GEN_1627; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1629 = 4'h7 == _T_89777 ? shiftedStoreDataQPreg_7 : _GEN_1628; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1630 = 4'h8 == _T_89777 ? shiftedStoreDataQPreg_8 : _GEN_1629; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1631 = 4'h9 == _T_89777 ? shiftedStoreDataQPreg_9 : _GEN_1630; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1632 = 4'ha == _T_89777 ? shiftedStoreDataQPreg_10 : _GEN_1631; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1633 = 4'hb == _T_89777 ? shiftedStoreDataQPreg_11 : _GEN_1632; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1634 = 4'hc == _T_89777 ? shiftedStoreDataQPreg_12 : _GEN_1633; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1635 = 4'hd == _T_89777 ? shiftedStoreDataQPreg_13 : _GEN_1634; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1636 = 4'he == _T_89777 ? shiftedStoreDataQPreg_14 : _GEN_1635; // @[LoadQueue.scala 195:31:@38771.6]
  assign _GEN_1637 = 4'hf == _T_89777 ? shiftedStoreDataQPreg_15 : _GEN_1636; // @[LoadQueue.scala 195:31:@38771.6]
  assign lastConflict_11_0 = _T_89794 ? _GEN_1590 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_1 = _T_89794 ? _GEN_1591 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_2 = _T_89794 ? _GEN_1592 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_3 = _T_89794 ? _GEN_1593 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_4 = _T_89794 ? _GEN_1594 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_5 = _T_89794 ? _GEN_1595 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_6 = _T_89794 ? _GEN_1596 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_7 = _T_89794 ? _GEN_1597 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_8 = _T_89794 ? _GEN_1598 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_9 = _T_89794 ? _GEN_1599 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_10 = _T_89794 ? _GEN_1600 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_11 = _T_89794 ? _GEN_1601 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_12 = _T_89794 ? _GEN_1602 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_13 = _T_89794 ? _GEN_1603 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_14 = _T_89794 ? _GEN_1604 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign lastConflict_11_15 = _T_89794 ? _GEN_1605 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign canBypass_11 = _T_89794 ? _GEN_1621 : 1'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign bypassVal_11 = _T_89794 ? _GEN_1637 : 32'h0; // @[LoadQueue.scala 192:53:@38768.4]
  assign _T_89900 = conflictPReg_12_2 ? 2'h2 : {{1'd0}, conflictPReg_12_1}; // @[LoadQueue.scala 191:60:@38825.4]
  assign _T_89901 = conflictPReg_12_3 ? 2'h3 : _T_89900; // @[LoadQueue.scala 191:60:@38826.4]
  assign _T_89902 = conflictPReg_12_4 ? 3'h4 : {{1'd0}, _T_89901}; // @[LoadQueue.scala 191:60:@38827.4]
  assign _T_89903 = conflictPReg_12_5 ? 3'h5 : _T_89902; // @[LoadQueue.scala 191:60:@38828.4]
  assign _T_89904 = conflictPReg_12_6 ? 3'h6 : _T_89903; // @[LoadQueue.scala 191:60:@38829.4]
  assign _T_89905 = conflictPReg_12_7 ? 3'h7 : _T_89904; // @[LoadQueue.scala 191:60:@38830.4]
  assign _T_89906 = conflictPReg_12_8 ? 4'h8 : {{1'd0}, _T_89905}; // @[LoadQueue.scala 191:60:@38831.4]
  assign _T_89907 = conflictPReg_12_9 ? 4'h9 : _T_89906; // @[LoadQueue.scala 191:60:@38832.4]
  assign _T_89908 = conflictPReg_12_10 ? 4'ha : _T_89907; // @[LoadQueue.scala 191:60:@38833.4]
  assign _T_89909 = conflictPReg_12_11 ? 4'hb : _T_89908; // @[LoadQueue.scala 191:60:@38834.4]
  assign _T_89910 = conflictPReg_12_12 ? 4'hc : _T_89909; // @[LoadQueue.scala 191:60:@38835.4]
  assign _T_89911 = conflictPReg_12_13 ? 4'hd : _T_89910; // @[LoadQueue.scala 191:60:@38836.4]
  assign _T_89912 = conflictPReg_12_14 ? 4'he : _T_89911; // @[LoadQueue.scala 191:60:@38837.4]
  assign _T_89913 = conflictPReg_12_15 ? 4'hf : _T_89912; // @[LoadQueue.scala 191:60:@38838.4]
  assign _T_89916 = conflictPReg_12_0 | conflictPReg_12_1; // @[LoadQueue.scala 192:43:@38840.4]
  assign _T_89917 = _T_89916 | conflictPReg_12_2; // @[LoadQueue.scala 192:43:@38841.4]
  assign _T_89918 = _T_89917 | conflictPReg_12_3; // @[LoadQueue.scala 192:43:@38842.4]
  assign _T_89919 = _T_89918 | conflictPReg_12_4; // @[LoadQueue.scala 192:43:@38843.4]
  assign _T_89920 = _T_89919 | conflictPReg_12_5; // @[LoadQueue.scala 192:43:@38844.4]
  assign _T_89921 = _T_89920 | conflictPReg_12_6; // @[LoadQueue.scala 192:43:@38845.4]
  assign _T_89922 = _T_89921 | conflictPReg_12_7; // @[LoadQueue.scala 192:43:@38846.4]
  assign _T_89923 = _T_89922 | conflictPReg_12_8; // @[LoadQueue.scala 192:43:@38847.4]
  assign _T_89924 = _T_89923 | conflictPReg_12_9; // @[LoadQueue.scala 192:43:@38848.4]
  assign _T_89925 = _T_89924 | conflictPReg_12_10; // @[LoadQueue.scala 192:43:@38849.4]
  assign _T_89926 = _T_89925 | conflictPReg_12_11; // @[LoadQueue.scala 192:43:@38850.4]
  assign _T_89927 = _T_89926 | conflictPReg_12_12; // @[LoadQueue.scala 192:43:@38851.4]
  assign _T_89928 = _T_89927 | conflictPReg_12_13; // @[LoadQueue.scala 192:43:@38852.4]
  assign _T_89929 = _T_89928 | conflictPReg_12_14; // @[LoadQueue.scala 192:43:@38853.4]
  assign _T_89930 = _T_89929 | conflictPReg_12_15; // @[LoadQueue.scala 192:43:@38854.4]
  assign _GEN_1656 = 4'h0 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1657 = 4'h1 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1658 = 4'h2 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1659 = 4'h3 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1660 = 4'h4 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1661 = 4'h5 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1662 = 4'h6 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1663 = 4'h7 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1664 = 4'h8 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1665 = 4'h9 == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1666 = 4'ha == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1667 = 4'hb == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1668 = 4'hc == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1669 = 4'hd == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1670 = 4'he == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1671 = 4'hf == _T_89913; // @[LoadQueue.scala 193:43:@38856.6]
  assign _GEN_1673 = 4'h1 == _T_89913 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1674 = 4'h2 == _T_89913 ? shiftedStoreDataKnownPReg_2 : _GEN_1673; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1675 = 4'h3 == _T_89913 ? shiftedStoreDataKnownPReg_3 : _GEN_1674; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1676 = 4'h4 == _T_89913 ? shiftedStoreDataKnownPReg_4 : _GEN_1675; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1677 = 4'h5 == _T_89913 ? shiftedStoreDataKnownPReg_5 : _GEN_1676; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1678 = 4'h6 == _T_89913 ? shiftedStoreDataKnownPReg_6 : _GEN_1677; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1679 = 4'h7 == _T_89913 ? shiftedStoreDataKnownPReg_7 : _GEN_1678; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1680 = 4'h8 == _T_89913 ? shiftedStoreDataKnownPReg_8 : _GEN_1679; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1681 = 4'h9 == _T_89913 ? shiftedStoreDataKnownPReg_9 : _GEN_1680; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1682 = 4'ha == _T_89913 ? shiftedStoreDataKnownPReg_10 : _GEN_1681; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1683 = 4'hb == _T_89913 ? shiftedStoreDataKnownPReg_11 : _GEN_1682; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1684 = 4'hc == _T_89913 ? shiftedStoreDataKnownPReg_12 : _GEN_1683; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1685 = 4'hd == _T_89913 ? shiftedStoreDataKnownPReg_13 : _GEN_1684; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1686 = 4'he == _T_89913 ? shiftedStoreDataKnownPReg_14 : _GEN_1685; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1687 = 4'hf == _T_89913 ? shiftedStoreDataKnownPReg_15 : _GEN_1686; // @[LoadQueue.scala 194:31:@38857.6]
  assign _GEN_1689 = 4'h1 == _T_89913 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1690 = 4'h2 == _T_89913 ? shiftedStoreDataQPreg_2 : _GEN_1689; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1691 = 4'h3 == _T_89913 ? shiftedStoreDataQPreg_3 : _GEN_1690; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1692 = 4'h4 == _T_89913 ? shiftedStoreDataQPreg_4 : _GEN_1691; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1693 = 4'h5 == _T_89913 ? shiftedStoreDataQPreg_5 : _GEN_1692; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1694 = 4'h6 == _T_89913 ? shiftedStoreDataQPreg_6 : _GEN_1693; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1695 = 4'h7 == _T_89913 ? shiftedStoreDataQPreg_7 : _GEN_1694; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1696 = 4'h8 == _T_89913 ? shiftedStoreDataQPreg_8 : _GEN_1695; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1697 = 4'h9 == _T_89913 ? shiftedStoreDataQPreg_9 : _GEN_1696; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1698 = 4'ha == _T_89913 ? shiftedStoreDataQPreg_10 : _GEN_1697; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1699 = 4'hb == _T_89913 ? shiftedStoreDataQPreg_11 : _GEN_1698; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1700 = 4'hc == _T_89913 ? shiftedStoreDataQPreg_12 : _GEN_1699; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1701 = 4'hd == _T_89913 ? shiftedStoreDataQPreg_13 : _GEN_1700; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1702 = 4'he == _T_89913 ? shiftedStoreDataQPreg_14 : _GEN_1701; // @[LoadQueue.scala 195:31:@38858.6]
  assign _GEN_1703 = 4'hf == _T_89913 ? shiftedStoreDataQPreg_15 : _GEN_1702; // @[LoadQueue.scala 195:31:@38858.6]
  assign lastConflict_12_0 = _T_89930 ? _GEN_1656 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_1 = _T_89930 ? _GEN_1657 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_2 = _T_89930 ? _GEN_1658 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_3 = _T_89930 ? _GEN_1659 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_4 = _T_89930 ? _GEN_1660 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_5 = _T_89930 ? _GEN_1661 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_6 = _T_89930 ? _GEN_1662 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_7 = _T_89930 ? _GEN_1663 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_8 = _T_89930 ? _GEN_1664 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_9 = _T_89930 ? _GEN_1665 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_10 = _T_89930 ? _GEN_1666 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_11 = _T_89930 ? _GEN_1667 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_12 = _T_89930 ? _GEN_1668 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_13 = _T_89930 ? _GEN_1669 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_14 = _T_89930 ? _GEN_1670 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign lastConflict_12_15 = _T_89930 ? _GEN_1671 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign canBypass_12 = _T_89930 ? _GEN_1687 : 1'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign bypassVal_12 = _T_89930 ? _GEN_1703 : 32'h0; // @[LoadQueue.scala 192:53:@38855.4]
  assign _T_90036 = conflictPReg_13_2 ? 2'h2 : {{1'd0}, conflictPReg_13_1}; // @[LoadQueue.scala 191:60:@38912.4]
  assign _T_90037 = conflictPReg_13_3 ? 2'h3 : _T_90036; // @[LoadQueue.scala 191:60:@38913.4]
  assign _T_90038 = conflictPReg_13_4 ? 3'h4 : {{1'd0}, _T_90037}; // @[LoadQueue.scala 191:60:@38914.4]
  assign _T_90039 = conflictPReg_13_5 ? 3'h5 : _T_90038; // @[LoadQueue.scala 191:60:@38915.4]
  assign _T_90040 = conflictPReg_13_6 ? 3'h6 : _T_90039; // @[LoadQueue.scala 191:60:@38916.4]
  assign _T_90041 = conflictPReg_13_7 ? 3'h7 : _T_90040; // @[LoadQueue.scala 191:60:@38917.4]
  assign _T_90042 = conflictPReg_13_8 ? 4'h8 : {{1'd0}, _T_90041}; // @[LoadQueue.scala 191:60:@38918.4]
  assign _T_90043 = conflictPReg_13_9 ? 4'h9 : _T_90042; // @[LoadQueue.scala 191:60:@38919.4]
  assign _T_90044 = conflictPReg_13_10 ? 4'ha : _T_90043; // @[LoadQueue.scala 191:60:@38920.4]
  assign _T_90045 = conflictPReg_13_11 ? 4'hb : _T_90044; // @[LoadQueue.scala 191:60:@38921.4]
  assign _T_90046 = conflictPReg_13_12 ? 4'hc : _T_90045; // @[LoadQueue.scala 191:60:@38922.4]
  assign _T_90047 = conflictPReg_13_13 ? 4'hd : _T_90046; // @[LoadQueue.scala 191:60:@38923.4]
  assign _T_90048 = conflictPReg_13_14 ? 4'he : _T_90047; // @[LoadQueue.scala 191:60:@38924.4]
  assign _T_90049 = conflictPReg_13_15 ? 4'hf : _T_90048; // @[LoadQueue.scala 191:60:@38925.4]
  assign _T_90052 = conflictPReg_13_0 | conflictPReg_13_1; // @[LoadQueue.scala 192:43:@38927.4]
  assign _T_90053 = _T_90052 | conflictPReg_13_2; // @[LoadQueue.scala 192:43:@38928.4]
  assign _T_90054 = _T_90053 | conflictPReg_13_3; // @[LoadQueue.scala 192:43:@38929.4]
  assign _T_90055 = _T_90054 | conflictPReg_13_4; // @[LoadQueue.scala 192:43:@38930.4]
  assign _T_90056 = _T_90055 | conflictPReg_13_5; // @[LoadQueue.scala 192:43:@38931.4]
  assign _T_90057 = _T_90056 | conflictPReg_13_6; // @[LoadQueue.scala 192:43:@38932.4]
  assign _T_90058 = _T_90057 | conflictPReg_13_7; // @[LoadQueue.scala 192:43:@38933.4]
  assign _T_90059 = _T_90058 | conflictPReg_13_8; // @[LoadQueue.scala 192:43:@38934.4]
  assign _T_90060 = _T_90059 | conflictPReg_13_9; // @[LoadQueue.scala 192:43:@38935.4]
  assign _T_90061 = _T_90060 | conflictPReg_13_10; // @[LoadQueue.scala 192:43:@38936.4]
  assign _T_90062 = _T_90061 | conflictPReg_13_11; // @[LoadQueue.scala 192:43:@38937.4]
  assign _T_90063 = _T_90062 | conflictPReg_13_12; // @[LoadQueue.scala 192:43:@38938.4]
  assign _T_90064 = _T_90063 | conflictPReg_13_13; // @[LoadQueue.scala 192:43:@38939.4]
  assign _T_90065 = _T_90064 | conflictPReg_13_14; // @[LoadQueue.scala 192:43:@38940.4]
  assign _T_90066 = _T_90065 | conflictPReg_13_15; // @[LoadQueue.scala 192:43:@38941.4]
  assign _GEN_1722 = 4'h0 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1723 = 4'h1 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1724 = 4'h2 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1725 = 4'h3 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1726 = 4'h4 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1727 = 4'h5 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1728 = 4'h6 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1729 = 4'h7 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1730 = 4'h8 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1731 = 4'h9 == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1732 = 4'ha == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1733 = 4'hb == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1734 = 4'hc == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1735 = 4'hd == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1736 = 4'he == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1737 = 4'hf == _T_90049; // @[LoadQueue.scala 193:43:@38943.6]
  assign _GEN_1739 = 4'h1 == _T_90049 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1740 = 4'h2 == _T_90049 ? shiftedStoreDataKnownPReg_2 : _GEN_1739; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1741 = 4'h3 == _T_90049 ? shiftedStoreDataKnownPReg_3 : _GEN_1740; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1742 = 4'h4 == _T_90049 ? shiftedStoreDataKnownPReg_4 : _GEN_1741; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1743 = 4'h5 == _T_90049 ? shiftedStoreDataKnownPReg_5 : _GEN_1742; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1744 = 4'h6 == _T_90049 ? shiftedStoreDataKnownPReg_6 : _GEN_1743; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1745 = 4'h7 == _T_90049 ? shiftedStoreDataKnownPReg_7 : _GEN_1744; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1746 = 4'h8 == _T_90049 ? shiftedStoreDataKnownPReg_8 : _GEN_1745; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1747 = 4'h9 == _T_90049 ? shiftedStoreDataKnownPReg_9 : _GEN_1746; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1748 = 4'ha == _T_90049 ? shiftedStoreDataKnownPReg_10 : _GEN_1747; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1749 = 4'hb == _T_90049 ? shiftedStoreDataKnownPReg_11 : _GEN_1748; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1750 = 4'hc == _T_90049 ? shiftedStoreDataKnownPReg_12 : _GEN_1749; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1751 = 4'hd == _T_90049 ? shiftedStoreDataKnownPReg_13 : _GEN_1750; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1752 = 4'he == _T_90049 ? shiftedStoreDataKnownPReg_14 : _GEN_1751; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1753 = 4'hf == _T_90049 ? shiftedStoreDataKnownPReg_15 : _GEN_1752; // @[LoadQueue.scala 194:31:@38944.6]
  assign _GEN_1755 = 4'h1 == _T_90049 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1756 = 4'h2 == _T_90049 ? shiftedStoreDataQPreg_2 : _GEN_1755; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1757 = 4'h3 == _T_90049 ? shiftedStoreDataQPreg_3 : _GEN_1756; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1758 = 4'h4 == _T_90049 ? shiftedStoreDataQPreg_4 : _GEN_1757; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1759 = 4'h5 == _T_90049 ? shiftedStoreDataQPreg_5 : _GEN_1758; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1760 = 4'h6 == _T_90049 ? shiftedStoreDataQPreg_6 : _GEN_1759; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1761 = 4'h7 == _T_90049 ? shiftedStoreDataQPreg_7 : _GEN_1760; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1762 = 4'h8 == _T_90049 ? shiftedStoreDataQPreg_8 : _GEN_1761; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1763 = 4'h9 == _T_90049 ? shiftedStoreDataQPreg_9 : _GEN_1762; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1764 = 4'ha == _T_90049 ? shiftedStoreDataQPreg_10 : _GEN_1763; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1765 = 4'hb == _T_90049 ? shiftedStoreDataQPreg_11 : _GEN_1764; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1766 = 4'hc == _T_90049 ? shiftedStoreDataQPreg_12 : _GEN_1765; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1767 = 4'hd == _T_90049 ? shiftedStoreDataQPreg_13 : _GEN_1766; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1768 = 4'he == _T_90049 ? shiftedStoreDataQPreg_14 : _GEN_1767; // @[LoadQueue.scala 195:31:@38945.6]
  assign _GEN_1769 = 4'hf == _T_90049 ? shiftedStoreDataQPreg_15 : _GEN_1768; // @[LoadQueue.scala 195:31:@38945.6]
  assign lastConflict_13_0 = _T_90066 ? _GEN_1722 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_1 = _T_90066 ? _GEN_1723 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_2 = _T_90066 ? _GEN_1724 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_3 = _T_90066 ? _GEN_1725 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_4 = _T_90066 ? _GEN_1726 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_5 = _T_90066 ? _GEN_1727 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_6 = _T_90066 ? _GEN_1728 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_7 = _T_90066 ? _GEN_1729 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_8 = _T_90066 ? _GEN_1730 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_9 = _T_90066 ? _GEN_1731 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_10 = _T_90066 ? _GEN_1732 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_11 = _T_90066 ? _GEN_1733 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_12 = _T_90066 ? _GEN_1734 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_13 = _T_90066 ? _GEN_1735 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_14 = _T_90066 ? _GEN_1736 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign lastConflict_13_15 = _T_90066 ? _GEN_1737 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign canBypass_13 = _T_90066 ? _GEN_1753 : 1'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign bypassVal_13 = _T_90066 ? _GEN_1769 : 32'h0; // @[LoadQueue.scala 192:53:@38942.4]
  assign _T_90172 = conflictPReg_14_2 ? 2'h2 : {{1'd0}, conflictPReg_14_1}; // @[LoadQueue.scala 191:60:@38999.4]
  assign _T_90173 = conflictPReg_14_3 ? 2'h3 : _T_90172; // @[LoadQueue.scala 191:60:@39000.4]
  assign _T_90174 = conflictPReg_14_4 ? 3'h4 : {{1'd0}, _T_90173}; // @[LoadQueue.scala 191:60:@39001.4]
  assign _T_90175 = conflictPReg_14_5 ? 3'h5 : _T_90174; // @[LoadQueue.scala 191:60:@39002.4]
  assign _T_90176 = conflictPReg_14_6 ? 3'h6 : _T_90175; // @[LoadQueue.scala 191:60:@39003.4]
  assign _T_90177 = conflictPReg_14_7 ? 3'h7 : _T_90176; // @[LoadQueue.scala 191:60:@39004.4]
  assign _T_90178 = conflictPReg_14_8 ? 4'h8 : {{1'd0}, _T_90177}; // @[LoadQueue.scala 191:60:@39005.4]
  assign _T_90179 = conflictPReg_14_9 ? 4'h9 : _T_90178; // @[LoadQueue.scala 191:60:@39006.4]
  assign _T_90180 = conflictPReg_14_10 ? 4'ha : _T_90179; // @[LoadQueue.scala 191:60:@39007.4]
  assign _T_90181 = conflictPReg_14_11 ? 4'hb : _T_90180; // @[LoadQueue.scala 191:60:@39008.4]
  assign _T_90182 = conflictPReg_14_12 ? 4'hc : _T_90181; // @[LoadQueue.scala 191:60:@39009.4]
  assign _T_90183 = conflictPReg_14_13 ? 4'hd : _T_90182; // @[LoadQueue.scala 191:60:@39010.4]
  assign _T_90184 = conflictPReg_14_14 ? 4'he : _T_90183; // @[LoadQueue.scala 191:60:@39011.4]
  assign _T_90185 = conflictPReg_14_15 ? 4'hf : _T_90184; // @[LoadQueue.scala 191:60:@39012.4]
  assign _T_90188 = conflictPReg_14_0 | conflictPReg_14_1; // @[LoadQueue.scala 192:43:@39014.4]
  assign _T_90189 = _T_90188 | conflictPReg_14_2; // @[LoadQueue.scala 192:43:@39015.4]
  assign _T_90190 = _T_90189 | conflictPReg_14_3; // @[LoadQueue.scala 192:43:@39016.4]
  assign _T_90191 = _T_90190 | conflictPReg_14_4; // @[LoadQueue.scala 192:43:@39017.4]
  assign _T_90192 = _T_90191 | conflictPReg_14_5; // @[LoadQueue.scala 192:43:@39018.4]
  assign _T_90193 = _T_90192 | conflictPReg_14_6; // @[LoadQueue.scala 192:43:@39019.4]
  assign _T_90194 = _T_90193 | conflictPReg_14_7; // @[LoadQueue.scala 192:43:@39020.4]
  assign _T_90195 = _T_90194 | conflictPReg_14_8; // @[LoadQueue.scala 192:43:@39021.4]
  assign _T_90196 = _T_90195 | conflictPReg_14_9; // @[LoadQueue.scala 192:43:@39022.4]
  assign _T_90197 = _T_90196 | conflictPReg_14_10; // @[LoadQueue.scala 192:43:@39023.4]
  assign _T_90198 = _T_90197 | conflictPReg_14_11; // @[LoadQueue.scala 192:43:@39024.4]
  assign _T_90199 = _T_90198 | conflictPReg_14_12; // @[LoadQueue.scala 192:43:@39025.4]
  assign _T_90200 = _T_90199 | conflictPReg_14_13; // @[LoadQueue.scala 192:43:@39026.4]
  assign _T_90201 = _T_90200 | conflictPReg_14_14; // @[LoadQueue.scala 192:43:@39027.4]
  assign _T_90202 = _T_90201 | conflictPReg_14_15; // @[LoadQueue.scala 192:43:@39028.4]
  assign _GEN_1788 = 4'h0 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1789 = 4'h1 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1790 = 4'h2 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1791 = 4'h3 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1792 = 4'h4 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1793 = 4'h5 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1794 = 4'h6 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1795 = 4'h7 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1796 = 4'h8 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1797 = 4'h9 == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1798 = 4'ha == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1799 = 4'hb == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1800 = 4'hc == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1801 = 4'hd == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1802 = 4'he == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1803 = 4'hf == _T_90185; // @[LoadQueue.scala 193:43:@39030.6]
  assign _GEN_1805 = 4'h1 == _T_90185 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1806 = 4'h2 == _T_90185 ? shiftedStoreDataKnownPReg_2 : _GEN_1805; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1807 = 4'h3 == _T_90185 ? shiftedStoreDataKnownPReg_3 : _GEN_1806; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1808 = 4'h4 == _T_90185 ? shiftedStoreDataKnownPReg_4 : _GEN_1807; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1809 = 4'h5 == _T_90185 ? shiftedStoreDataKnownPReg_5 : _GEN_1808; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1810 = 4'h6 == _T_90185 ? shiftedStoreDataKnownPReg_6 : _GEN_1809; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1811 = 4'h7 == _T_90185 ? shiftedStoreDataKnownPReg_7 : _GEN_1810; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1812 = 4'h8 == _T_90185 ? shiftedStoreDataKnownPReg_8 : _GEN_1811; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1813 = 4'h9 == _T_90185 ? shiftedStoreDataKnownPReg_9 : _GEN_1812; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1814 = 4'ha == _T_90185 ? shiftedStoreDataKnownPReg_10 : _GEN_1813; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1815 = 4'hb == _T_90185 ? shiftedStoreDataKnownPReg_11 : _GEN_1814; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1816 = 4'hc == _T_90185 ? shiftedStoreDataKnownPReg_12 : _GEN_1815; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1817 = 4'hd == _T_90185 ? shiftedStoreDataKnownPReg_13 : _GEN_1816; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1818 = 4'he == _T_90185 ? shiftedStoreDataKnownPReg_14 : _GEN_1817; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1819 = 4'hf == _T_90185 ? shiftedStoreDataKnownPReg_15 : _GEN_1818; // @[LoadQueue.scala 194:31:@39031.6]
  assign _GEN_1821 = 4'h1 == _T_90185 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1822 = 4'h2 == _T_90185 ? shiftedStoreDataQPreg_2 : _GEN_1821; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1823 = 4'h3 == _T_90185 ? shiftedStoreDataQPreg_3 : _GEN_1822; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1824 = 4'h4 == _T_90185 ? shiftedStoreDataQPreg_4 : _GEN_1823; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1825 = 4'h5 == _T_90185 ? shiftedStoreDataQPreg_5 : _GEN_1824; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1826 = 4'h6 == _T_90185 ? shiftedStoreDataQPreg_6 : _GEN_1825; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1827 = 4'h7 == _T_90185 ? shiftedStoreDataQPreg_7 : _GEN_1826; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1828 = 4'h8 == _T_90185 ? shiftedStoreDataQPreg_8 : _GEN_1827; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1829 = 4'h9 == _T_90185 ? shiftedStoreDataQPreg_9 : _GEN_1828; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1830 = 4'ha == _T_90185 ? shiftedStoreDataQPreg_10 : _GEN_1829; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1831 = 4'hb == _T_90185 ? shiftedStoreDataQPreg_11 : _GEN_1830; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1832 = 4'hc == _T_90185 ? shiftedStoreDataQPreg_12 : _GEN_1831; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1833 = 4'hd == _T_90185 ? shiftedStoreDataQPreg_13 : _GEN_1832; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1834 = 4'he == _T_90185 ? shiftedStoreDataQPreg_14 : _GEN_1833; // @[LoadQueue.scala 195:31:@39032.6]
  assign _GEN_1835 = 4'hf == _T_90185 ? shiftedStoreDataQPreg_15 : _GEN_1834; // @[LoadQueue.scala 195:31:@39032.6]
  assign lastConflict_14_0 = _T_90202 ? _GEN_1788 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_1 = _T_90202 ? _GEN_1789 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_2 = _T_90202 ? _GEN_1790 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_3 = _T_90202 ? _GEN_1791 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_4 = _T_90202 ? _GEN_1792 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_5 = _T_90202 ? _GEN_1793 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_6 = _T_90202 ? _GEN_1794 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_7 = _T_90202 ? _GEN_1795 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_8 = _T_90202 ? _GEN_1796 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_9 = _T_90202 ? _GEN_1797 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_10 = _T_90202 ? _GEN_1798 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_11 = _T_90202 ? _GEN_1799 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_12 = _T_90202 ? _GEN_1800 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_13 = _T_90202 ? _GEN_1801 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_14 = _T_90202 ? _GEN_1802 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign lastConflict_14_15 = _T_90202 ? _GEN_1803 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign canBypass_14 = _T_90202 ? _GEN_1819 : 1'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign bypassVal_14 = _T_90202 ? _GEN_1835 : 32'h0; // @[LoadQueue.scala 192:53:@39029.4]
  assign _T_90308 = conflictPReg_15_2 ? 2'h2 : {{1'd0}, conflictPReg_15_1}; // @[LoadQueue.scala 191:60:@39086.4]
  assign _T_90309 = conflictPReg_15_3 ? 2'h3 : _T_90308; // @[LoadQueue.scala 191:60:@39087.4]
  assign _T_90310 = conflictPReg_15_4 ? 3'h4 : {{1'd0}, _T_90309}; // @[LoadQueue.scala 191:60:@39088.4]
  assign _T_90311 = conflictPReg_15_5 ? 3'h5 : _T_90310; // @[LoadQueue.scala 191:60:@39089.4]
  assign _T_90312 = conflictPReg_15_6 ? 3'h6 : _T_90311; // @[LoadQueue.scala 191:60:@39090.4]
  assign _T_90313 = conflictPReg_15_7 ? 3'h7 : _T_90312; // @[LoadQueue.scala 191:60:@39091.4]
  assign _T_90314 = conflictPReg_15_8 ? 4'h8 : {{1'd0}, _T_90313}; // @[LoadQueue.scala 191:60:@39092.4]
  assign _T_90315 = conflictPReg_15_9 ? 4'h9 : _T_90314; // @[LoadQueue.scala 191:60:@39093.4]
  assign _T_90316 = conflictPReg_15_10 ? 4'ha : _T_90315; // @[LoadQueue.scala 191:60:@39094.4]
  assign _T_90317 = conflictPReg_15_11 ? 4'hb : _T_90316; // @[LoadQueue.scala 191:60:@39095.4]
  assign _T_90318 = conflictPReg_15_12 ? 4'hc : _T_90317; // @[LoadQueue.scala 191:60:@39096.4]
  assign _T_90319 = conflictPReg_15_13 ? 4'hd : _T_90318; // @[LoadQueue.scala 191:60:@39097.4]
  assign _T_90320 = conflictPReg_15_14 ? 4'he : _T_90319; // @[LoadQueue.scala 191:60:@39098.4]
  assign _T_90321 = conflictPReg_15_15 ? 4'hf : _T_90320; // @[LoadQueue.scala 191:60:@39099.4]
  assign _T_90324 = conflictPReg_15_0 | conflictPReg_15_1; // @[LoadQueue.scala 192:43:@39101.4]
  assign _T_90325 = _T_90324 | conflictPReg_15_2; // @[LoadQueue.scala 192:43:@39102.4]
  assign _T_90326 = _T_90325 | conflictPReg_15_3; // @[LoadQueue.scala 192:43:@39103.4]
  assign _T_90327 = _T_90326 | conflictPReg_15_4; // @[LoadQueue.scala 192:43:@39104.4]
  assign _T_90328 = _T_90327 | conflictPReg_15_5; // @[LoadQueue.scala 192:43:@39105.4]
  assign _T_90329 = _T_90328 | conflictPReg_15_6; // @[LoadQueue.scala 192:43:@39106.4]
  assign _T_90330 = _T_90329 | conflictPReg_15_7; // @[LoadQueue.scala 192:43:@39107.4]
  assign _T_90331 = _T_90330 | conflictPReg_15_8; // @[LoadQueue.scala 192:43:@39108.4]
  assign _T_90332 = _T_90331 | conflictPReg_15_9; // @[LoadQueue.scala 192:43:@39109.4]
  assign _T_90333 = _T_90332 | conflictPReg_15_10; // @[LoadQueue.scala 192:43:@39110.4]
  assign _T_90334 = _T_90333 | conflictPReg_15_11; // @[LoadQueue.scala 192:43:@39111.4]
  assign _T_90335 = _T_90334 | conflictPReg_15_12; // @[LoadQueue.scala 192:43:@39112.4]
  assign _T_90336 = _T_90335 | conflictPReg_15_13; // @[LoadQueue.scala 192:43:@39113.4]
  assign _T_90337 = _T_90336 | conflictPReg_15_14; // @[LoadQueue.scala 192:43:@39114.4]
  assign _T_90338 = _T_90337 | conflictPReg_15_15; // @[LoadQueue.scala 192:43:@39115.4]
  assign _GEN_1854 = 4'h0 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1855 = 4'h1 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1856 = 4'h2 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1857 = 4'h3 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1858 = 4'h4 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1859 = 4'h5 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1860 = 4'h6 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1861 = 4'h7 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1862 = 4'h8 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1863 = 4'h9 == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1864 = 4'ha == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1865 = 4'hb == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1866 = 4'hc == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1867 = 4'hd == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1868 = 4'he == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1869 = 4'hf == _T_90321; // @[LoadQueue.scala 193:43:@39117.6]
  assign _GEN_1871 = 4'h1 == _T_90321 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1872 = 4'h2 == _T_90321 ? shiftedStoreDataKnownPReg_2 : _GEN_1871; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1873 = 4'h3 == _T_90321 ? shiftedStoreDataKnownPReg_3 : _GEN_1872; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1874 = 4'h4 == _T_90321 ? shiftedStoreDataKnownPReg_4 : _GEN_1873; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1875 = 4'h5 == _T_90321 ? shiftedStoreDataKnownPReg_5 : _GEN_1874; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1876 = 4'h6 == _T_90321 ? shiftedStoreDataKnownPReg_6 : _GEN_1875; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1877 = 4'h7 == _T_90321 ? shiftedStoreDataKnownPReg_7 : _GEN_1876; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1878 = 4'h8 == _T_90321 ? shiftedStoreDataKnownPReg_8 : _GEN_1877; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1879 = 4'h9 == _T_90321 ? shiftedStoreDataKnownPReg_9 : _GEN_1878; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1880 = 4'ha == _T_90321 ? shiftedStoreDataKnownPReg_10 : _GEN_1879; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1881 = 4'hb == _T_90321 ? shiftedStoreDataKnownPReg_11 : _GEN_1880; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1882 = 4'hc == _T_90321 ? shiftedStoreDataKnownPReg_12 : _GEN_1881; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1883 = 4'hd == _T_90321 ? shiftedStoreDataKnownPReg_13 : _GEN_1882; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1884 = 4'he == _T_90321 ? shiftedStoreDataKnownPReg_14 : _GEN_1883; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1885 = 4'hf == _T_90321 ? shiftedStoreDataKnownPReg_15 : _GEN_1884; // @[LoadQueue.scala 194:31:@39118.6]
  assign _GEN_1887 = 4'h1 == _T_90321 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1888 = 4'h2 == _T_90321 ? shiftedStoreDataQPreg_2 : _GEN_1887; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1889 = 4'h3 == _T_90321 ? shiftedStoreDataQPreg_3 : _GEN_1888; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1890 = 4'h4 == _T_90321 ? shiftedStoreDataQPreg_4 : _GEN_1889; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1891 = 4'h5 == _T_90321 ? shiftedStoreDataQPreg_5 : _GEN_1890; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1892 = 4'h6 == _T_90321 ? shiftedStoreDataQPreg_6 : _GEN_1891; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1893 = 4'h7 == _T_90321 ? shiftedStoreDataQPreg_7 : _GEN_1892; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1894 = 4'h8 == _T_90321 ? shiftedStoreDataQPreg_8 : _GEN_1893; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1895 = 4'h9 == _T_90321 ? shiftedStoreDataQPreg_9 : _GEN_1894; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1896 = 4'ha == _T_90321 ? shiftedStoreDataQPreg_10 : _GEN_1895; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1897 = 4'hb == _T_90321 ? shiftedStoreDataQPreg_11 : _GEN_1896; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1898 = 4'hc == _T_90321 ? shiftedStoreDataQPreg_12 : _GEN_1897; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1899 = 4'hd == _T_90321 ? shiftedStoreDataQPreg_13 : _GEN_1898; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1900 = 4'he == _T_90321 ? shiftedStoreDataQPreg_14 : _GEN_1899; // @[LoadQueue.scala 195:31:@39119.6]
  assign _GEN_1901 = 4'hf == _T_90321 ? shiftedStoreDataQPreg_15 : _GEN_1900; // @[LoadQueue.scala 195:31:@39119.6]
  assign lastConflict_15_0 = _T_90338 ? _GEN_1854 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_1 = _T_90338 ? _GEN_1855 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_2 = _T_90338 ? _GEN_1856 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_3 = _T_90338 ? _GEN_1857 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_4 = _T_90338 ? _GEN_1858 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_5 = _T_90338 ? _GEN_1859 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_6 = _T_90338 ? _GEN_1860 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_7 = _T_90338 ? _GEN_1861 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_8 = _T_90338 ? _GEN_1862 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_9 = _T_90338 ? _GEN_1863 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_10 = _T_90338 ? _GEN_1864 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_11 = _T_90338 ? _GEN_1865 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_12 = _T_90338 ? _GEN_1866 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_13 = _T_90338 ? _GEN_1867 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_14 = _T_90338 ? _GEN_1868 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign lastConflict_15_15 = _T_90338 ? _GEN_1869 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign canBypass_15 = _T_90338 ? _GEN_1885 : 1'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign bypassVal_15 = _T_90338 ? _GEN_1901 : 32'h0; // @[LoadQueue.scala 192:53:@39116.4]
  assign _T_90398 = 16'h1 << head; // @[OneHot.scala 52:12:@39124.4]
  assign _T_90400 = _T_90398[0]; // @[util.scala 33:60:@39126.4]
  assign _T_90401 = _T_90398[1]; // @[util.scala 33:60:@39127.4]
  assign _T_90402 = _T_90398[2]; // @[util.scala 33:60:@39128.4]
  assign _T_90403 = _T_90398[3]; // @[util.scala 33:60:@39129.4]
  assign _T_90404 = _T_90398[4]; // @[util.scala 33:60:@39130.4]
  assign _T_90405 = _T_90398[5]; // @[util.scala 33:60:@39131.4]
  assign _T_90406 = _T_90398[6]; // @[util.scala 33:60:@39132.4]
  assign _T_90407 = _T_90398[7]; // @[util.scala 33:60:@39133.4]
  assign _T_90408 = _T_90398[8]; // @[util.scala 33:60:@39134.4]
  assign _T_90409 = _T_90398[9]; // @[util.scala 33:60:@39135.4]
  assign _T_90410 = _T_90398[10]; // @[util.scala 33:60:@39136.4]
  assign _T_90411 = _T_90398[11]; // @[util.scala 33:60:@39137.4]
  assign _T_90412 = _T_90398[12]; // @[util.scala 33:60:@39138.4]
  assign _T_90413 = _T_90398[13]; // @[util.scala 33:60:@39139.4]
  assign _T_90414 = _T_90398[14]; // @[util.scala 33:60:@39140.4]
  assign _T_90415 = _T_90398[15]; // @[util.scala 33:60:@39141.4]
  assign _T_93512 = dataKnownPReg_15 == 1'h0; // @[LoadQueue.scala 229:41:@41664.4]
  assign _T_93513 = addrKnownPReg_15 & _T_93512; // @[LoadQueue.scala 229:38:@41665.4]
  assign _T_93515 = bypassInitiated_15 == 1'h0; // @[LoadQueue.scala 230:12:@41667.6]
  assign _T_93517 = prevPriorityRequest_15 == 1'h0; // @[LoadQueue.scala 230:46:@41668.6]
  assign _T_93518 = _T_93515 & _T_93517; // @[LoadQueue.scala 230:43:@41669.6]
  assign _T_93520 = dataKnown_15 == 1'h0; // @[LoadQueue.scala 230:84:@41670.6]
  assign _T_93521 = _T_93518 & _T_93520; // @[LoadQueue.scala 230:81:@41671.6]
  assign _T_93524 = storeAddrNotKnownFlagsPReg_15_0 | storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 233:86:@41674.8]
  assign _T_93525 = _T_93524 | storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 233:86:@41675.8]
  assign _T_93526 = _T_93525 | storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 233:86:@41676.8]
  assign _T_93527 = _T_93526 | storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 233:86:@41677.8]
  assign _T_93528 = _T_93527 | storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 233:86:@41678.8]
  assign _T_93529 = _T_93528 | storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 233:86:@41679.8]
  assign _T_93530 = _T_93529 | storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 233:86:@41680.8]
  assign _T_93531 = _T_93530 | storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 233:86:@41681.8]
  assign _T_93532 = _T_93531 | storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 233:86:@41682.8]
  assign _T_93533 = _T_93532 | storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 233:86:@41683.8]
  assign _T_93534 = _T_93533 | storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 233:86:@41684.8]
  assign _T_93535 = _T_93534 | storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 233:86:@41685.8]
  assign _T_93536 = _T_93535 | storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 233:86:@41686.8]
  assign _T_93537 = _T_93536 | storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 233:86:@41687.8]
  assign _T_93538 = _T_93537 | storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 233:86:@41688.8]
  assign _T_93540 = _T_93538 == 1'h0; // @[LoadQueue.scala 233:38:@41689.8]
  assign _T_93559 = _T_90338 == 1'h0; // @[LoadQueue.scala 234:11:@41706.8]
  assign _T_93560 = _T_93540 & _T_93559; // @[LoadQueue.scala 233:103:@41707.8]
  assign _GEN_2028 = _T_93521 ? _T_93560 : 1'h0; // @[LoadQueue.scala 230:110:@41672.6]
  assign loadRequest_15 = _T_93513 ? _GEN_2028 : 1'h0; // @[LoadQueue.scala 229:71:@41666.4]
  assign _T_90456 = loadRequest_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39159.4]
  assign _T_93428 = dataKnownPReg_14 == 1'h0; // @[LoadQueue.scala 229:41:@41582.4]
  assign _T_93429 = addrKnownPReg_14 & _T_93428; // @[LoadQueue.scala 229:38:@41583.4]
  assign _T_93431 = bypassInitiated_14 == 1'h0; // @[LoadQueue.scala 230:12:@41585.6]
  assign _T_93433 = prevPriorityRequest_14 == 1'h0; // @[LoadQueue.scala 230:46:@41586.6]
  assign _T_93434 = _T_93431 & _T_93433; // @[LoadQueue.scala 230:43:@41587.6]
  assign _T_93436 = dataKnown_14 == 1'h0; // @[LoadQueue.scala 230:84:@41588.6]
  assign _T_93437 = _T_93434 & _T_93436; // @[LoadQueue.scala 230:81:@41589.6]
  assign _T_93440 = storeAddrNotKnownFlagsPReg_14_0 | storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 233:86:@41592.8]
  assign _T_93441 = _T_93440 | storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 233:86:@41593.8]
  assign _T_93442 = _T_93441 | storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 233:86:@41594.8]
  assign _T_93443 = _T_93442 | storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 233:86:@41595.8]
  assign _T_93444 = _T_93443 | storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 233:86:@41596.8]
  assign _T_93445 = _T_93444 | storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 233:86:@41597.8]
  assign _T_93446 = _T_93445 | storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 233:86:@41598.8]
  assign _T_93447 = _T_93446 | storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 233:86:@41599.8]
  assign _T_93448 = _T_93447 | storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 233:86:@41600.8]
  assign _T_93449 = _T_93448 | storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 233:86:@41601.8]
  assign _T_93450 = _T_93449 | storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 233:86:@41602.8]
  assign _T_93451 = _T_93450 | storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 233:86:@41603.8]
  assign _T_93452 = _T_93451 | storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 233:86:@41604.8]
  assign _T_93453 = _T_93452 | storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 233:86:@41605.8]
  assign _T_93454 = _T_93453 | storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 233:86:@41606.8]
  assign _T_93456 = _T_93454 == 1'h0; // @[LoadQueue.scala 233:38:@41607.8]
  assign _T_93475 = _T_90202 == 1'h0; // @[LoadQueue.scala 234:11:@41624.8]
  assign _T_93476 = _T_93456 & _T_93475; // @[LoadQueue.scala 233:103:@41625.8]
  assign _GEN_2024 = _T_93437 ? _T_93476 : 1'h0; // @[LoadQueue.scala 230:110:@41590.6]
  assign loadRequest_14 = _T_93429 ? _GEN_2024 : 1'h0; // @[LoadQueue.scala 229:71:@41584.4]
  assign _T_90457 = loadRequest_14 ? 16'h4000 : _T_90456; // @[Mux.scala 31:69:@39160.4]
  assign _T_93344 = dataKnownPReg_13 == 1'h0; // @[LoadQueue.scala 229:41:@41500.4]
  assign _T_93345 = addrKnownPReg_13 & _T_93344; // @[LoadQueue.scala 229:38:@41501.4]
  assign _T_93347 = bypassInitiated_13 == 1'h0; // @[LoadQueue.scala 230:12:@41503.6]
  assign _T_93349 = prevPriorityRequest_13 == 1'h0; // @[LoadQueue.scala 230:46:@41504.6]
  assign _T_93350 = _T_93347 & _T_93349; // @[LoadQueue.scala 230:43:@41505.6]
  assign _T_93352 = dataKnown_13 == 1'h0; // @[LoadQueue.scala 230:84:@41506.6]
  assign _T_93353 = _T_93350 & _T_93352; // @[LoadQueue.scala 230:81:@41507.6]
  assign _T_93356 = storeAddrNotKnownFlagsPReg_13_0 | storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 233:86:@41510.8]
  assign _T_93357 = _T_93356 | storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 233:86:@41511.8]
  assign _T_93358 = _T_93357 | storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 233:86:@41512.8]
  assign _T_93359 = _T_93358 | storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 233:86:@41513.8]
  assign _T_93360 = _T_93359 | storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 233:86:@41514.8]
  assign _T_93361 = _T_93360 | storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 233:86:@41515.8]
  assign _T_93362 = _T_93361 | storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 233:86:@41516.8]
  assign _T_93363 = _T_93362 | storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 233:86:@41517.8]
  assign _T_93364 = _T_93363 | storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 233:86:@41518.8]
  assign _T_93365 = _T_93364 | storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 233:86:@41519.8]
  assign _T_93366 = _T_93365 | storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 233:86:@41520.8]
  assign _T_93367 = _T_93366 | storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 233:86:@41521.8]
  assign _T_93368 = _T_93367 | storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 233:86:@41522.8]
  assign _T_93369 = _T_93368 | storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 233:86:@41523.8]
  assign _T_93370 = _T_93369 | storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 233:86:@41524.8]
  assign _T_93372 = _T_93370 == 1'h0; // @[LoadQueue.scala 233:38:@41525.8]
  assign _T_93391 = _T_90066 == 1'h0; // @[LoadQueue.scala 234:11:@41542.8]
  assign _T_93392 = _T_93372 & _T_93391; // @[LoadQueue.scala 233:103:@41543.8]
  assign _GEN_2020 = _T_93353 ? _T_93392 : 1'h0; // @[LoadQueue.scala 230:110:@41508.6]
  assign loadRequest_13 = _T_93345 ? _GEN_2020 : 1'h0; // @[LoadQueue.scala 229:71:@41502.4]
  assign _T_90458 = loadRequest_13 ? 16'h2000 : _T_90457; // @[Mux.scala 31:69:@39161.4]
  assign _T_93260 = dataKnownPReg_12 == 1'h0; // @[LoadQueue.scala 229:41:@41418.4]
  assign _T_93261 = addrKnownPReg_12 & _T_93260; // @[LoadQueue.scala 229:38:@41419.4]
  assign _T_93263 = bypassInitiated_12 == 1'h0; // @[LoadQueue.scala 230:12:@41421.6]
  assign _T_93265 = prevPriorityRequest_12 == 1'h0; // @[LoadQueue.scala 230:46:@41422.6]
  assign _T_93266 = _T_93263 & _T_93265; // @[LoadQueue.scala 230:43:@41423.6]
  assign _T_93268 = dataKnown_12 == 1'h0; // @[LoadQueue.scala 230:84:@41424.6]
  assign _T_93269 = _T_93266 & _T_93268; // @[LoadQueue.scala 230:81:@41425.6]
  assign _T_93272 = storeAddrNotKnownFlagsPReg_12_0 | storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 233:86:@41428.8]
  assign _T_93273 = _T_93272 | storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 233:86:@41429.8]
  assign _T_93274 = _T_93273 | storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 233:86:@41430.8]
  assign _T_93275 = _T_93274 | storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 233:86:@41431.8]
  assign _T_93276 = _T_93275 | storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 233:86:@41432.8]
  assign _T_93277 = _T_93276 | storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 233:86:@41433.8]
  assign _T_93278 = _T_93277 | storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 233:86:@41434.8]
  assign _T_93279 = _T_93278 | storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 233:86:@41435.8]
  assign _T_93280 = _T_93279 | storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 233:86:@41436.8]
  assign _T_93281 = _T_93280 | storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 233:86:@41437.8]
  assign _T_93282 = _T_93281 | storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 233:86:@41438.8]
  assign _T_93283 = _T_93282 | storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 233:86:@41439.8]
  assign _T_93284 = _T_93283 | storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 233:86:@41440.8]
  assign _T_93285 = _T_93284 | storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 233:86:@41441.8]
  assign _T_93286 = _T_93285 | storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 233:86:@41442.8]
  assign _T_93288 = _T_93286 == 1'h0; // @[LoadQueue.scala 233:38:@41443.8]
  assign _T_93307 = _T_89930 == 1'h0; // @[LoadQueue.scala 234:11:@41460.8]
  assign _T_93308 = _T_93288 & _T_93307; // @[LoadQueue.scala 233:103:@41461.8]
  assign _GEN_2016 = _T_93269 ? _T_93308 : 1'h0; // @[LoadQueue.scala 230:110:@41426.6]
  assign loadRequest_12 = _T_93261 ? _GEN_2016 : 1'h0; // @[LoadQueue.scala 229:71:@41420.4]
  assign _T_90459 = loadRequest_12 ? 16'h1000 : _T_90458; // @[Mux.scala 31:69:@39162.4]
  assign _T_93176 = dataKnownPReg_11 == 1'h0; // @[LoadQueue.scala 229:41:@41336.4]
  assign _T_93177 = addrKnownPReg_11 & _T_93176; // @[LoadQueue.scala 229:38:@41337.4]
  assign _T_93179 = bypassInitiated_11 == 1'h0; // @[LoadQueue.scala 230:12:@41339.6]
  assign _T_93181 = prevPriorityRequest_11 == 1'h0; // @[LoadQueue.scala 230:46:@41340.6]
  assign _T_93182 = _T_93179 & _T_93181; // @[LoadQueue.scala 230:43:@41341.6]
  assign _T_93184 = dataKnown_11 == 1'h0; // @[LoadQueue.scala 230:84:@41342.6]
  assign _T_93185 = _T_93182 & _T_93184; // @[LoadQueue.scala 230:81:@41343.6]
  assign _T_93188 = storeAddrNotKnownFlagsPReg_11_0 | storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 233:86:@41346.8]
  assign _T_93189 = _T_93188 | storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 233:86:@41347.8]
  assign _T_93190 = _T_93189 | storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 233:86:@41348.8]
  assign _T_93191 = _T_93190 | storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 233:86:@41349.8]
  assign _T_93192 = _T_93191 | storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 233:86:@41350.8]
  assign _T_93193 = _T_93192 | storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 233:86:@41351.8]
  assign _T_93194 = _T_93193 | storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 233:86:@41352.8]
  assign _T_93195 = _T_93194 | storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 233:86:@41353.8]
  assign _T_93196 = _T_93195 | storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 233:86:@41354.8]
  assign _T_93197 = _T_93196 | storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 233:86:@41355.8]
  assign _T_93198 = _T_93197 | storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 233:86:@41356.8]
  assign _T_93199 = _T_93198 | storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 233:86:@41357.8]
  assign _T_93200 = _T_93199 | storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 233:86:@41358.8]
  assign _T_93201 = _T_93200 | storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 233:86:@41359.8]
  assign _T_93202 = _T_93201 | storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 233:86:@41360.8]
  assign _T_93204 = _T_93202 == 1'h0; // @[LoadQueue.scala 233:38:@41361.8]
  assign _T_93223 = _T_89794 == 1'h0; // @[LoadQueue.scala 234:11:@41378.8]
  assign _T_93224 = _T_93204 & _T_93223; // @[LoadQueue.scala 233:103:@41379.8]
  assign _GEN_2012 = _T_93185 ? _T_93224 : 1'h0; // @[LoadQueue.scala 230:110:@41344.6]
  assign loadRequest_11 = _T_93177 ? _GEN_2012 : 1'h0; // @[LoadQueue.scala 229:71:@41338.4]
  assign _T_90460 = loadRequest_11 ? 16'h800 : _T_90459; // @[Mux.scala 31:69:@39163.4]
  assign _T_93092 = dataKnownPReg_10 == 1'h0; // @[LoadQueue.scala 229:41:@41254.4]
  assign _T_93093 = addrKnownPReg_10 & _T_93092; // @[LoadQueue.scala 229:38:@41255.4]
  assign _T_93095 = bypassInitiated_10 == 1'h0; // @[LoadQueue.scala 230:12:@41257.6]
  assign _T_93097 = prevPriorityRequest_10 == 1'h0; // @[LoadQueue.scala 230:46:@41258.6]
  assign _T_93098 = _T_93095 & _T_93097; // @[LoadQueue.scala 230:43:@41259.6]
  assign _T_93100 = dataKnown_10 == 1'h0; // @[LoadQueue.scala 230:84:@41260.6]
  assign _T_93101 = _T_93098 & _T_93100; // @[LoadQueue.scala 230:81:@41261.6]
  assign _T_93104 = storeAddrNotKnownFlagsPReg_10_0 | storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 233:86:@41264.8]
  assign _T_93105 = _T_93104 | storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 233:86:@41265.8]
  assign _T_93106 = _T_93105 | storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 233:86:@41266.8]
  assign _T_93107 = _T_93106 | storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 233:86:@41267.8]
  assign _T_93108 = _T_93107 | storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 233:86:@41268.8]
  assign _T_93109 = _T_93108 | storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 233:86:@41269.8]
  assign _T_93110 = _T_93109 | storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 233:86:@41270.8]
  assign _T_93111 = _T_93110 | storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 233:86:@41271.8]
  assign _T_93112 = _T_93111 | storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 233:86:@41272.8]
  assign _T_93113 = _T_93112 | storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 233:86:@41273.8]
  assign _T_93114 = _T_93113 | storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 233:86:@41274.8]
  assign _T_93115 = _T_93114 | storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 233:86:@41275.8]
  assign _T_93116 = _T_93115 | storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 233:86:@41276.8]
  assign _T_93117 = _T_93116 | storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 233:86:@41277.8]
  assign _T_93118 = _T_93117 | storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 233:86:@41278.8]
  assign _T_93120 = _T_93118 == 1'h0; // @[LoadQueue.scala 233:38:@41279.8]
  assign _T_93139 = _T_89658 == 1'h0; // @[LoadQueue.scala 234:11:@41296.8]
  assign _T_93140 = _T_93120 & _T_93139; // @[LoadQueue.scala 233:103:@41297.8]
  assign _GEN_2008 = _T_93101 ? _T_93140 : 1'h0; // @[LoadQueue.scala 230:110:@41262.6]
  assign loadRequest_10 = _T_93093 ? _GEN_2008 : 1'h0; // @[LoadQueue.scala 229:71:@41256.4]
  assign _T_90461 = loadRequest_10 ? 16'h400 : _T_90460; // @[Mux.scala 31:69:@39164.4]
  assign _T_93008 = dataKnownPReg_9 == 1'h0; // @[LoadQueue.scala 229:41:@41172.4]
  assign _T_93009 = addrKnownPReg_9 & _T_93008; // @[LoadQueue.scala 229:38:@41173.4]
  assign _T_93011 = bypassInitiated_9 == 1'h0; // @[LoadQueue.scala 230:12:@41175.6]
  assign _T_93013 = prevPriorityRequest_9 == 1'h0; // @[LoadQueue.scala 230:46:@41176.6]
  assign _T_93014 = _T_93011 & _T_93013; // @[LoadQueue.scala 230:43:@41177.6]
  assign _T_93016 = dataKnown_9 == 1'h0; // @[LoadQueue.scala 230:84:@41178.6]
  assign _T_93017 = _T_93014 & _T_93016; // @[LoadQueue.scala 230:81:@41179.6]
  assign _T_93020 = storeAddrNotKnownFlagsPReg_9_0 | storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 233:86:@41182.8]
  assign _T_93021 = _T_93020 | storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 233:86:@41183.8]
  assign _T_93022 = _T_93021 | storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 233:86:@41184.8]
  assign _T_93023 = _T_93022 | storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 233:86:@41185.8]
  assign _T_93024 = _T_93023 | storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 233:86:@41186.8]
  assign _T_93025 = _T_93024 | storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 233:86:@41187.8]
  assign _T_93026 = _T_93025 | storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 233:86:@41188.8]
  assign _T_93027 = _T_93026 | storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 233:86:@41189.8]
  assign _T_93028 = _T_93027 | storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 233:86:@41190.8]
  assign _T_93029 = _T_93028 | storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 233:86:@41191.8]
  assign _T_93030 = _T_93029 | storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 233:86:@41192.8]
  assign _T_93031 = _T_93030 | storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 233:86:@41193.8]
  assign _T_93032 = _T_93031 | storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 233:86:@41194.8]
  assign _T_93033 = _T_93032 | storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 233:86:@41195.8]
  assign _T_93034 = _T_93033 | storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 233:86:@41196.8]
  assign _T_93036 = _T_93034 == 1'h0; // @[LoadQueue.scala 233:38:@41197.8]
  assign _T_93055 = _T_89522 == 1'h0; // @[LoadQueue.scala 234:11:@41214.8]
  assign _T_93056 = _T_93036 & _T_93055; // @[LoadQueue.scala 233:103:@41215.8]
  assign _GEN_2004 = _T_93017 ? _T_93056 : 1'h0; // @[LoadQueue.scala 230:110:@41180.6]
  assign loadRequest_9 = _T_93009 ? _GEN_2004 : 1'h0; // @[LoadQueue.scala 229:71:@41174.4]
  assign _T_90462 = loadRequest_9 ? 16'h200 : _T_90461; // @[Mux.scala 31:69:@39165.4]
  assign _T_92924 = dataKnownPReg_8 == 1'h0; // @[LoadQueue.scala 229:41:@41090.4]
  assign _T_92925 = addrKnownPReg_8 & _T_92924; // @[LoadQueue.scala 229:38:@41091.4]
  assign _T_92927 = bypassInitiated_8 == 1'h0; // @[LoadQueue.scala 230:12:@41093.6]
  assign _T_92929 = prevPriorityRequest_8 == 1'h0; // @[LoadQueue.scala 230:46:@41094.6]
  assign _T_92930 = _T_92927 & _T_92929; // @[LoadQueue.scala 230:43:@41095.6]
  assign _T_92932 = dataKnown_8 == 1'h0; // @[LoadQueue.scala 230:84:@41096.6]
  assign _T_92933 = _T_92930 & _T_92932; // @[LoadQueue.scala 230:81:@41097.6]
  assign _T_92936 = storeAddrNotKnownFlagsPReg_8_0 | storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 233:86:@41100.8]
  assign _T_92937 = _T_92936 | storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 233:86:@41101.8]
  assign _T_92938 = _T_92937 | storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 233:86:@41102.8]
  assign _T_92939 = _T_92938 | storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 233:86:@41103.8]
  assign _T_92940 = _T_92939 | storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 233:86:@41104.8]
  assign _T_92941 = _T_92940 | storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 233:86:@41105.8]
  assign _T_92942 = _T_92941 | storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 233:86:@41106.8]
  assign _T_92943 = _T_92942 | storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 233:86:@41107.8]
  assign _T_92944 = _T_92943 | storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 233:86:@41108.8]
  assign _T_92945 = _T_92944 | storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 233:86:@41109.8]
  assign _T_92946 = _T_92945 | storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 233:86:@41110.8]
  assign _T_92947 = _T_92946 | storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 233:86:@41111.8]
  assign _T_92948 = _T_92947 | storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 233:86:@41112.8]
  assign _T_92949 = _T_92948 | storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 233:86:@41113.8]
  assign _T_92950 = _T_92949 | storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 233:86:@41114.8]
  assign _T_92952 = _T_92950 == 1'h0; // @[LoadQueue.scala 233:38:@41115.8]
  assign _T_92971 = _T_89386 == 1'h0; // @[LoadQueue.scala 234:11:@41132.8]
  assign _T_92972 = _T_92952 & _T_92971; // @[LoadQueue.scala 233:103:@41133.8]
  assign _GEN_2000 = _T_92933 ? _T_92972 : 1'h0; // @[LoadQueue.scala 230:110:@41098.6]
  assign loadRequest_8 = _T_92925 ? _GEN_2000 : 1'h0; // @[LoadQueue.scala 229:71:@41092.4]
  assign _T_90463 = loadRequest_8 ? 16'h100 : _T_90462; // @[Mux.scala 31:69:@39166.4]
  assign _T_92840 = dataKnownPReg_7 == 1'h0; // @[LoadQueue.scala 229:41:@41008.4]
  assign _T_92841 = addrKnownPReg_7 & _T_92840; // @[LoadQueue.scala 229:38:@41009.4]
  assign _T_92843 = bypassInitiated_7 == 1'h0; // @[LoadQueue.scala 230:12:@41011.6]
  assign _T_92845 = prevPriorityRequest_7 == 1'h0; // @[LoadQueue.scala 230:46:@41012.6]
  assign _T_92846 = _T_92843 & _T_92845; // @[LoadQueue.scala 230:43:@41013.6]
  assign _T_92848 = dataKnown_7 == 1'h0; // @[LoadQueue.scala 230:84:@41014.6]
  assign _T_92849 = _T_92846 & _T_92848; // @[LoadQueue.scala 230:81:@41015.6]
  assign _T_92852 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 233:86:@41018.8]
  assign _T_92853 = _T_92852 | storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 233:86:@41019.8]
  assign _T_92854 = _T_92853 | storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 233:86:@41020.8]
  assign _T_92855 = _T_92854 | storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 233:86:@41021.8]
  assign _T_92856 = _T_92855 | storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 233:86:@41022.8]
  assign _T_92857 = _T_92856 | storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 233:86:@41023.8]
  assign _T_92858 = _T_92857 | storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 233:86:@41024.8]
  assign _T_92859 = _T_92858 | storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 233:86:@41025.8]
  assign _T_92860 = _T_92859 | storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 233:86:@41026.8]
  assign _T_92861 = _T_92860 | storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 233:86:@41027.8]
  assign _T_92862 = _T_92861 | storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 233:86:@41028.8]
  assign _T_92863 = _T_92862 | storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 233:86:@41029.8]
  assign _T_92864 = _T_92863 | storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 233:86:@41030.8]
  assign _T_92865 = _T_92864 | storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 233:86:@41031.8]
  assign _T_92866 = _T_92865 | storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 233:86:@41032.8]
  assign _T_92868 = _T_92866 == 1'h0; // @[LoadQueue.scala 233:38:@41033.8]
  assign _T_92887 = _T_89250 == 1'h0; // @[LoadQueue.scala 234:11:@41050.8]
  assign _T_92888 = _T_92868 & _T_92887; // @[LoadQueue.scala 233:103:@41051.8]
  assign _GEN_1996 = _T_92849 ? _T_92888 : 1'h0; // @[LoadQueue.scala 230:110:@41016.6]
  assign loadRequest_7 = _T_92841 ? _GEN_1996 : 1'h0; // @[LoadQueue.scala 229:71:@41010.4]
  assign _T_90464 = loadRequest_7 ? 16'h80 : _T_90463; // @[Mux.scala 31:69:@39167.4]
  assign _T_92756 = dataKnownPReg_6 == 1'h0; // @[LoadQueue.scala 229:41:@40926.4]
  assign _T_92757 = addrKnownPReg_6 & _T_92756; // @[LoadQueue.scala 229:38:@40927.4]
  assign _T_92759 = bypassInitiated_6 == 1'h0; // @[LoadQueue.scala 230:12:@40929.6]
  assign _T_92761 = prevPriorityRequest_6 == 1'h0; // @[LoadQueue.scala 230:46:@40930.6]
  assign _T_92762 = _T_92759 & _T_92761; // @[LoadQueue.scala 230:43:@40931.6]
  assign _T_92764 = dataKnown_6 == 1'h0; // @[LoadQueue.scala 230:84:@40932.6]
  assign _T_92765 = _T_92762 & _T_92764; // @[LoadQueue.scala 230:81:@40933.6]
  assign _T_92768 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 233:86:@40936.8]
  assign _T_92769 = _T_92768 | storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 233:86:@40937.8]
  assign _T_92770 = _T_92769 | storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 233:86:@40938.8]
  assign _T_92771 = _T_92770 | storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 233:86:@40939.8]
  assign _T_92772 = _T_92771 | storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 233:86:@40940.8]
  assign _T_92773 = _T_92772 | storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 233:86:@40941.8]
  assign _T_92774 = _T_92773 | storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 233:86:@40942.8]
  assign _T_92775 = _T_92774 | storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 233:86:@40943.8]
  assign _T_92776 = _T_92775 | storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 233:86:@40944.8]
  assign _T_92777 = _T_92776 | storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 233:86:@40945.8]
  assign _T_92778 = _T_92777 | storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 233:86:@40946.8]
  assign _T_92779 = _T_92778 | storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 233:86:@40947.8]
  assign _T_92780 = _T_92779 | storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 233:86:@40948.8]
  assign _T_92781 = _T_92780 | storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 233:86:@40949.8]
  assign _T_92782 = _T_92781 | storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 233:86:@40950.8]
  assign _T_92784 = _T_92782 == 1'h0; // @[LoadQueue.scala 233:38:@40951.8]
  assign _T_92803 = _T_89114 == 1'h0; // @[LoadQueue.scala 234:11:@40968.8]
  assign _T_92804 = _T_92784 & _T_92803; // @[LoadQueue.scala 233:103:@40969.8]
  assign _GEN_1992 = _T_92765 ? _T_92804 : 1'h0; // @[LoadQueue.scala 230:110:@40934.6]
  assign loadRequest_6 = _T_92757 ? _GEN_1992 : 1'h0; // @[LoadQueue.scala 229:71:@40928.4]
  assign _T_90465 = loadRequest_6 ? 16'h40 : _T_90464; // @[Mux.scala 31:69:@39168.4]
  assign _T_92672 = dataKnownPReg_5 == 1'h0; // @[LoadQueue.scala 229:41:@40844.4]
  assign _T_92673 = addrKnownPReg_5 & _T_92672; // @[LoadQueue.scala 229:38:@40845.4]
  assign _T_92675 = bypassInitiated_5 == 1'h0; // @[LoadQueue.scala 230:12:@40847.6]
  assign _T_92677 = prevPriorityRequest_5 == 1'h0; // @[LoadQueue.scala 230:46:@40848.6]
  assign _T_92678 = _T_92675 & _T_92677; // @[LoadQueue.scala 230:43:@40849.6]
  assign _T_92680 = dataKnown_5 == 1'h0; // @[LoadQueue.scala 230:84:@40850.6]
  assign _T_92681 = _T_92678 & _T_92680; // @[LoadQueue.scala 230:81:@40851.6]
  assign _T_92684 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 233:86:@40854.8]
  assign _T_92685 = _T_92684 | storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 233:86:@40855.8]
  assign _T_92686 = _T_92685 | storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 233:86:@40856.8]
  assign _T_92687 = _T_92686 | storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 233:86:@40857.8]
  assign _T_92688 = _T_92687 | storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 233:86:@40858.8]
  assign _T_92689 = _T_92688 | storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 233:86:@40859.8]
  assign _T_92690 = _T_92689 | storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 233:86:@40860.8]
  assign _T_92691 = _T_92690 | storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 233:86:@40861.8]
  assign _T_92692 = _T_92691 | storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 233:86:@40862.8]
  assign _T_92693 = _T_92692 | storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 233:86:@40863.8]
  assign _T_92694 = _T_92693 | storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 233:86:@40864.8]
  assign _T_92695 = _T_92694 | storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 233:86:@40865.8]
  assign _T_92696 = _T_92695 | storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 233:86:@40866.8]
  assign _T_92697 = _T_92696 | storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 233:86:@40867.8]
  assign _T_92698 = _T_92697 | storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 233:86:@40868.8]
  assign _T_92700 = _T_92698 == 1'h0; // @[LoadQueue.scala 233:38:@40869.8]
  assign _T_92719 = _T_88978 == 1'h0; // @[LoadQueue.scala 234:11:@40886.8]
  assign _T_92720 = _T_92700 & _T_92719; // @[LoadQueue.scala 233:103:@40887.8]
  assign _GEN_1988 = _T_92681 ? _T_92720 : 1'h0; // @[LoadQueue.scala 230:110:@40852.6]
  assign loadRequest_5 = _T_92673 ? _GEN_1988 : 1'h0; // @[LoadQueue.scala 229:71:@40846.4]
  assign _T_90466 = loadRequest_5 ? 16'h20 : _T_90465; // @[Mux.scala 31:69:@39169.4]
  assign _T_92588 = dataKnownPReg_4 == 1'h0; // @[LoadQueue.scala 229:41:@40762.4]
  assign _T_92589 = addrKnownPReg_4 & _T_92588; // @[LoadQueue.scala 229:38:@40763.4]
  assign _T_92591 = bypassInitiated_4 == 1'h0; // @[LoadQueue.scala 230:12:@40765.6]
  assign _T_92593 = prevPriorityRequest_4 == 1'h0; // @[LoadQueue.scala 230:46:@40766.6]
  assign _T_92594 = _T_92591 & _T_92593; // @[LoadQueue.scala 230:43:@40767.6]
  assign _T_92596 = dataKnown_4 == 1'h0; // @[LoadQueue.scala 230:84:@40768.6]
  assign _T_92597 = _T_92594 & _T_92596; // @[LoadQueue.scala 230:81:@40769.6]
  assign _T_92600 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 233:86:@40772.8]
  assign _T_92601 = _T_92600 | storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 233:86:@40773.8]
  assign _T_92602 = _T_92601 | storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 233:86:@40774.8]
  assign _T_92603 = _T_92602 | storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 233:86:@40775.8]
  assign _T_92604 = _T_92603 | storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 233:86:@40776.8]
  assign _T_92605 = _T_92604 | storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 233:86:@40777.8]
  assign _T_92606 = _T_92605 | storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 233:86:@40778.8]
  assign _T_92607 = _T_92606 | storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 233:86:@40779.8]
  assign _T_92608 = _T_92607 | storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 233:86:@40780.8]
  assign _T_92609 = _T_92608 | storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 233:86:@40781.8]
  assign _T_92610 = _T_92609 | storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 233:86:@40782.8]
  assign _T_92611 = _T_92610 | storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 233:86:@40783.8]
  assign _T_92612 = _T_92611 | storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 233:86:@40784.8]
  assign _T_92613 = _T_92612 | storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 233:86:@40785.8]
  assign _T_92614 = _T_92613 | storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 233:86:@40786.8]
  assign _T_92616 = _T_92614 == 1'h0; // @[LoadQueue.scala 233:38:@40787.8]
  assign _T_92635 = _T_88842 == 1'h0; // @[LoadQueue.scala 234:11:@40804.8]
  assign _T_92636 = _T_92616 & _T_92635; // @[LoadQueue.scala 233:103:@40805.8]
  assign _GEN_1984 = _T_92597 ? _T_92636 : 1'h0; // @[LoadQueue.scala 230:110:@40770.6]
  assign loadRequest_4 = _T_92589 ? _GEN_1984 : 1'h0; // @[LoadQueue.scala 229:71:@40764.4]
  assign _T_90467 = loadRequest_4 ? 16'h10 : _T_90466; // @[Mux.scala 31:69:@39170.4]
  assign _T_92504 = dataKnownPReg_3 == 1'h0; // @[LoadQueue.scala 229:41:@40680.4]
  assign _T_92505 = addrKnownPReg_3 & _T_92504; // @[LoadQueue.scala 229:38:@40681.4]
  assign _T_92507 = bypassInitiated_3 == 1'h0; // @[LoadQueue.scala 230:12:@40683.6]
  assign _T_92509 = prevPriorityRequest_3 == 1'h0; // @[LoadQueue.scala 230:46:@40684.6]
  assign _T_92510 = _T_92507 & _T_92509; // @[LoadQueue.scala 230:43:@40685.6]
  assign _T_92512 = dataKnown_3 == 1'h0; // @[LoadQueue.scala 230:84:@40686.6]
  assign _T_92513 = _T_92510 & _T_92512; // @[LoadQueue.scala 230:81:@40687.6]
  assign _T_92516 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 233:86:@40690.8]
  assign _T_92517 = _T_92516 | storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 233:86:@40691.8]
  assign _T_92518 = _T_92517 | storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 233:86:@40692.8]
  assign _T_92519 = _T_92518 | storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 233:86:@40693.8]
  assign _T_92520 = _T_92519 | storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 233:86:@40694.8]
  assign _T_92521 = _T_92520 | storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 233:86:@40695.8]
  assign _T_92522 = _T_92521 | storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 233:86:@40696.8]
  assign _T_92523 = _T_92522 | storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 233:86:@40697.8]
  assign _T_92524 = _T_92523 | storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 233:86:@40698.8]
  assign _T_92525 = _T_92524 | storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 233:86:@40699.8]
  assign _T_92526 = _T_92525 | storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 233:86:@40700.8]
  assign _T_92527 = _T_92526 | storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 233:86:@40701.8]
  assign _T_92528 = _T_92527 | storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 233:86:@40702.8]
  assign _T_92529 = _T_92528 | storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 233:86:@40703.8]
  assign _T_92530 = _T_92529 | storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 233:86:@40704.8]
  assign _T_92532 = _T_92530 == 1'h0; // @[LoadQueue.scala 233:38:@40705.8]
  assign _T_92551 = _T_88706 == 1'h0; // @[LoadQueue.scala 234:11:@40722.8]
  assign _T_92552 = _T_92532 & _T_92551; // @[LoadQueue.scala 233:103:@40723.8]
  assign _GEN_1980 = _T_92513 ? _T_92552 : 1'h0; // @[LoadQueue.scala 230:110:@40688.6]
  assign loadRequest_3 = _T_92505 ? _GEN_1980 : 1'h0; // @[LoadQueue.scala 229:71:@40682.4]
  assign _T_90468 = loadRequest_3 ? 16'h8 : _T_90467; // @[Mux.scala 31:69:@39171.4]
  assign _T_92420 = dataKnownPReg_2 == 1'h0; // @[LoadQueue.scala 229:41:@40598.4]
  assign _T_92421 = addrKnownPReg_2 & _T_92420; // @[LoadQueue.scala 229:38:@40599.4]
  assign _T_92423 = bypassInitiated_2 == 1'h0; // @[LoadQueue.scala 230:12:@40601.6]
  assign _T_92425 = prevPriorityRequest_2 == 1'h0; // @[LoadQueue.scala 230:46:@40602.6]
  assign _T_92426 = _T_92423 & _T_92425; // @[LoadQueue.scala 230:43:@40603.6]
  assign _T_92428 = dataKnown_2 == 1'h0; // @[LoadQueue.scala 230:84:@40604.6]
  assign _T_92429 = _T_92426 & _T_92428; // @[LoadQueue.scala 230:81:@40605.6]
  assign _T_92432 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 233:86:@40608.8]
  assign _T_92433 = _T_92432 | storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 233:86:@40609.8]
  assign _T_92434 = _T_92433 | storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 233:86:@40610.8]
  assign _T_92435 = _T_92434 | storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 233:86:@40611.8]
  assign _T_92436 = _T_92435 | storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 233:86:@40612.8]
  assign _T_92437 = _T_92436 | storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 233:86:@40613.8]
  assign _T_92438 = _T_92437 | storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 233:86:@40614.8]
  assign _T_92439 = _T_92438 | storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 233:86:@40615.8]
  assign _T_92440 = _T_92439 | storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 233:86:@40616.8]
  assign _T_92441 = _T_92440 | storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 233:86:@40617.8]
  assign _T_92442 = _T_92441 | storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 233:86:@40618.8]
  assign _T_92443 = _T_92442 | storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 233:86:@40619.8]
  assign _T_92444 = _T_92443 | storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 233:86:@40620.8]
  assign _T_92445 = _T_92444 | storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 233:86:@40621.8]
  assign _T_92446 = _T_92445 | storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 233:86:@40622.8]
  assign _T_92448 = _T_92446 == 1'h0; // @[LoadQueue.scala 233:38:@40623.8]
  assign _T_92467 = _T_88570 == 1'h0; // @[LoadQueue.scala 234:11:@40640.8]
  assign _T_92468 = _T_92448 & _T_92467; // @[LoadQueue.scala 233:103:@40641.8]
  assign _GEN_1976 = _T_92429 ? _T_92468 : 1'h0; // @[LoadQueue.scala 230:110:@40606.6]
  assign loadRequest_2 = _T_92421 ? _GEN_1976 : 1'h0; // @[LoadQueue.scala 229:71:@40600.4]
  assign _T_90469 = loadRequest_2 ? 16'h4 : _T_90468; // @[Mux.scala 31:69:@39172.4]
  assign _T_92336 = dataKnownPReg_1 == 1'h0; // @[LoadQueue.scala 229:41:@40516.4]
  assign _T_92337 = addrKnownPReg_1 & _T_92336; // @[LoadQueue.scala 229:38:@40517.4]
  assign _T_92339 = bypassInitiated_1 == 1'h0; // @[LoadQueue.scala 230:12:@40519.6]
  assign _T_92341 = prevPriorityRequest_1 == 1'h0; // @[LoadQueue.scala 230:46:@40520.6]
  assign _T_92342 = _T_92339 & _T_92341; // @[LoadQueue.scala 230:43:@40521.6]
  assign _T_92344 = dataKnown_1 == 1'h0; // @[LoadQueue.scala 230:84:@40522.6]
  assign _T_92345 = _T_92342 & _T_92344; // @[LoadQueue.scala 230:81:@40523.6]
  assign _T_92348 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 233:86:@40526.8]
  assign _T_92349 = _T_92348 | storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 233:86:@40527.8]
  assign _T_92350 = _T_92349 | storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 233:86:@40528.8]
  assign _T_92351 = _T_92350 | storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 233:86:@40529.8]
  assign _T_92352 = _T_92351 | storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 233:86:@40530.8]
  assign _T_92353 = _T_92352 | storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 233:86:@40531.8]
  assign _T_92354 = _T_92353 | storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 233:86:@40532.8]
  assign _T_92355 = _T_92354 | storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 233:86:@40533.8]
  assign _T_92356 = _T_92355 | storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 233:86:@40534.8]
  assign _T_92357 = _T_92356 | storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 233:86:@40535.8]
  assign _T_92358 = _T_92357 | storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 233:86:@40536.8]
  assign _T_92359 = _T_92358 | storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 233:86:@40537.8]
  assign _T_92360 = _T_92359 | storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 233:86:@40538.8]
  assign _T_92361 = _T_92360 | storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 233:86:@40539.8]
  assign _T_92362 = _T_92361 | storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 233:86:@40540.8]
  assign _T_92364 = _T_92362 == 1'h0; // @[LoadQueue.scala 233:38:@40541.8]
  assign _T_92383 = _T_88434 == 1'h0; // @[LoadQueue.scala 234:11:@40558.8]
  assign _T_92384 = _T_92364 & _T_92383; // @[LoadQueue.scala 233:103:@40559.8]
  assign _GEN_1972 = _T_92345 ? _T_92384 : 1'h0; // @[LoadQueue.scala 230:110:@40524.6]
  assign loadRequest_1 = _T_92337 ? _GEN_1972 : 1'h0; // @[LoadQueue.scala 229:71:@40518.4]
  assign _T_90470 = loadRequest_1 ? 16'h2 : _T_90469; // @[Mux.scala 31:69:@39173.4]
  assign _T_92252 = dataKnownPReg_0 == 1'h0; // @[LoadQueue.scala 229:41:@40434.4]
  assign _T_92253 = addrKnownPReg_0 & _T_92252; // @[LoadQueue.scala 229:38:@40435.4]
  assign _T_92255 = bypassInitiated_0 == 1'h0; // @[LoadQueue.scala 230:12:@40437.6]
  assign _T_92257 = prevPriorityRequest_0 == 1'h0; // @[LoadQueue.scala 230:46:@40438.6]
  assign _T_92258 = _T_92255 & _T_92257; // @[LoadQueue.scala 230:43:@40439.6]
  assign _T_92260 = dataKnown_0 == 1'h0; // @[LoadQueue.scala 230:84:@40440.6]
  assign _T_92261 = _T_92258 & _T_92260; // @[LoadQueue.scala 230:81:@40441.6]
  assign _T_92264 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 233:86:@40444.8]
  assign _T_92265 = _T_92264 | storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 233:86:@40445.8]
  assign _T_92266 = _T_92265 | storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 233:86:@40446.8]
  assign _T_92267 = _T_92266 | storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 233:86:@40447.8]
  assign _T_92268 = _T_92267 | storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 233:86:@40448.8]
  assign _T_92269 = _T_92268 | storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 233:86:@40449.8]
  assign _T_92270 = _T_92269 | storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 233:86:@40450.8]
  assign _T_92271 = _T_92270 | storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 233:86:@40451.8]
  assign _T_92272 = _T_92271 | storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 233:86:@40452.8]
  assign _T_92273 = _T_92272 | storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 233:86:@40453.8]
  assign _T_92274 = _T_92273 | storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 233:86:@40454.8]
  assign _T_92275 = _T_92274 | storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 233:86:@40455.8]
  assign _T_92276 = _T_92275 | storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 233:86:@40456.8]
  assign _T_92277 = _T_92276 | storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 233:86:@40457.8]
  assign _T_92278 = _T_92277 | storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 233:86:@40458.8]
  assign _T_92280 = _T_92278 == 1'h0; // @[LoadQueue.scala 233:38:@40459.8]
  assign _T_92299 = _T_88298 == 1'h0; // @[LoadQueue.scala 234:11:@40476.8]
  assign _T_92300 = _T_92280 & _T_92299; // @[LoadQueue.scala 233:103:@40477.8]
  assign _GEN_1968 = _T_92261 ? _T_92300 : 1'h0; // @[LoadQueue.scala 230:110:@40442.6]
  assign loadRequest_0 = _T_92253 ? _GEN_1968 : 1'h0; // @[LoadQueue.scala 229:71:@40436.4]
  assign _T_90471 = loadRequest_0 ? 16'h1 : _T_90470; // @[Mux.scala 31:69:@39174.4]
  assign _T_90472 = _T_90471[0]; // @[OneHot.scala 66:30:@39175.4]
  assign _T_90473 = _T_90471[1]; // @[OneHot.scala 66:30:@39176.4]
  assign _T_90474 = _T_90471[2]; // @[OneHot.scala 66:30:@39177.4]
  assign _T_90475 = _T_90471[3]; // @[OneHot.scala 66:30:@39178.4]
  assign _T_90476 = _T_90471[4]; // @[OneHot.scala 66:30:@39179.4]
  assign _T_90477 = _T_90471[5]; // @[OneHot.scala 66:30:@39180.4]
  assign _T_90478 = _T_90471[6]; // @[OneHot.scala 66:30:@39181.4]
  assign _T_90479 = _T_90471[7]; // @[OneHot.scala 66:30:@39182.4]
  assign _T_90480 = _T_90471[8]; // @[OneHot.scala 66:30:@39183.4]
  assign _T_90481 = _T_90471[9]; // @[OneHot.scala 66:30:@39184.4]
  assign _T_90482 = _T_90471[10]; // @[OneHot.scala 66:30:@39185.4]
  assign _T_90483 = _T_90471[11]; // @[OneHot.scala 66:30:@39186.4]
  assign _T_90484 = _T_90471[12]; // @[OneHot.scala 66:30:@39187.4]
  assign _T_90485 = _T_90471[13]; // @[OneHot.scala 66:30:@39188.4]
  assign _T_90486 = _T_90471[14]; // @[OneHot.scala 66:30:@39189.4]
  assign _T_90487 = _T_90471[15]; // @[OneHot.scala 66:30:@39190.4]
  assign _T_90528 = loadRequest_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39208.4]
  assign _T_90529 = loadRequest_15 ? 16'h4000 : _T_90528; // @[Mux.scala 31:69:@39209.4]
  assign _T_90530 = loadRequest_14 ? 16'h2000 : _T_90529; // @[Mux.scala 31:69:@39210.4]
  assign _T_90531 = loadRequest_13 ? 16'h1000 : _T_90530; // @[Mux.scala 31:69:@39211.4]
  assign _T_90532 = loadRequest_12 ? 16'h800 : _T_90531; // @[Mux.scala 31:69:@39212.4]
  assign _T_90533 = loadRequest_11 ? 16'h400 : _T_90532; // @[Mux.scala 31:69:@39213.4]
  assign _T_90534 = loadRequest_10 ? 16'h200 : _T_90533; // @[Mux.scala 31:69:@39214.4]
  assign _T_90535 = loadRequest_9 ? 16'h100 : _T_90534; // @[Mux.scala 31:69:@39215.4]
  assign _T_90536 = loadRequest_8 ? 16'h80 : _T_90535; // @[Mux.scala 31:69:@39216.4]
  assign _T_90537 = loadRequest_7 ? 16'h40 : _T_90536; // @[Mux.scala 31:69:@39217.4]
  assign _T_90538 = loadRequest_6 ? 16'h20 : _T_90537; // @[Mux.scala 31:69:@39218.4]
  assign _T_90539 = loadRequest_5 ? 16'h10 : _T_90538; // @[Mux.scala 31:69:@39219.4]
  assign _T_90540 = loadRequest_4 ? 16'h8 : _T_90539; // @[Mux.scala 31:69:@39220.4]
  assign _T_90541 = loadRequest_3 ? 16'h4 : _T_90540; // @[Mux.scala 31:69:@39221.4]
  assign _T_90542 = loadRequest_2 ? 16'h2 : _T_90541; // @[Mux.scala 31:69:@39222.4]
  assign _T_90543 = loadRequest_1 ? 16'h1 : _T_90542; // @[Mux.scala 31:69:@39223.4]
  assign _T_90544 = _T_90543[0]; // @[OneHot.scala 66:30:@39224.4]
  assign _T_90545 = _T_90543[1]; // @[OneHot.scala 66:30:@39225.4]
  assign _T_90546 = _T_90543[2]; // @[OneHot.scala 66:30:@39226.4]
  assign _T_90547 = _T_90543[3]; // @[OneHot.scala 66:30:@39227.4]
  assign _T_90548 = _T_90543[4]; // @[OneHot.scala 66:30:@39228.4]
  assign _T_90549 = _T_90543[5]; // @[OneHot.scala 66:30:@39229.4]
  assign _T_90550 = _T_90543[6]; // @[OneHot.scala 66:30:@39230.4]
  assign _T_90551 = _T_90543[7]; // @[OneHot.scala 66:30:@39231.4]
  assign _T_90552 = _T_90543[8]; // @[OneHot.scala 66:30:@39232.4]
  assign _T_90553 = _T_90543[9]; // @[OneHot.scala 66:30:@39233.4]
  assign _T_90554 = _T_90543[10]; // @[OneHot.scala 66:30:@39234.4]
  assign _T_90555 = _T_90543[11]; // @[OneHot.scala 66:30:@39235.4]
  assign _T_90556 = _T_90543[12]; // @[OneHot.scala 66:30:@39236.4]
  assign _T_90557 = _T_90543[13]; // @[OneHot.scala 66:30:@39237.4]
  assign _T_90558 = _T_90543[14]; // @[OneHot.scala 66:30:@39238.4]
  assign _T_90559 = _T_90543[15]; // @[OneHot.scala 66:30:@39239.4]
  assign _T_90600 = loadRequest_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39257.4]
  assign _T_90601 = loadRequest_0 ? 16'h4000 : _T_90600; // @[Mux.scala 31:69:@39258.4]
  assign _T_90602 = loadRequest_15 ? 16'h2000 : _T_90601; // @[Mux.scala 31:69:@39259.4]
  assign _T_90603 = loadRequest_14 ? 16'h1000 : _T_90602; // @[Mux.scala 31:69:@39260.4]
  assign _T_90604 = loadRequest_13 ? 16'h800 : _T_90603; // @[Mux.scala 31:69:@39261.4]
  assign _T_90605 = loadRequest_12 ? 16'h400 : _T_90604; // @[Mux.scala 31:69:@39262.4]
  assign _T_90606 = loadRequest_11 ? 16'h200 : _T_90605; // @[Mux.scala 31:69:@39263.4]
  assign _T_90607 = loadRequest_10 ? 16'h100 : _T_90606; // @[Mux.scala 31:69:@39264.4]
  assign _T_90608 = loadRequest_9 ? 16'h80 : _T_90607; // @[Mux.scala 31:69:@39265.4]
  assign _T_90609 = loadRequest_8 ? 16'h40 : _T_90608; // @[Mux.scala 31:69:@39266.4]
  assign _T_90610 = loadRequest_7 ? 16'h20 : _T_90609; // @[Mux.scala 31:69:@39267.4]
  assign _T_90611 = loadRequest_6 ? 16'h10 : _T_90610; // @[Mux.scala 31:69:@39268.4]
  assign _T_90612 = loadRequest_5 ? 16'h8 : _T_90611; // @[Mux.scala 31:69:@39269.4]
  assign _T_90613 = loadRequest_4 ? 16'h4 : _T_90612; // @[Mux.scala 31:69:@39270.4]
  assign _T_90614 = loadRequest_3 ? 16'h2 : _T_90613; // @[Mux.scala 31:69:@39271.4]
  assign _T_90615 = loadRequest_2 ? 16'h1 : _T_90614; // @[Mux.scala 31:69:@39272.4]
  assign _T_90616 = _T_90615[0]; // @[OneHot.scala 66:30:@39273.4]
  assign _T_90617 = _T_90615[1]; // @[OneHot.scala 66:30:@39274.4]
  assign _T_90618 = _T_90615[2]; // @[OneHot.scala 66:30:@39275.4]
  assign _T_90619 = _T_90615[3]; // @[OneHot.scala 66:30:@39276.4]
  assign _T_90620 = _T_90615[4]; // @[OneHot.scala 66:30:@39277.4]
  assign _T_90621 = _T_90615[5]; // @[OneHot.scala 66:30:@39278.4]
  assign _T_90622 = _T_90615[6]; // @[OneHot.scala 66:30:@39279.4]
  assign _T_90623 = _T_90615[7]; // @[OneHot.scala 66:30:@39280.4]
  assign _T_90624 = _T_90615[8]; // @[OneHot.scala 66:30:@39281.4]
  assign _T_90625 = _T_90615[9]; // @[OneHot.scala 66:30:@39282.4]
  assign _T_90626 = _T_90615[10]; // @[OneHot.scala 66:30:@39283.4]
  assign _T_90627 = _T_90615[11]; // @[OneHot.scala 66:30:@39284.4]
  assign _T_90628 = _T_90615[12]; // @[OneHot.scala 66:30:@39285.4]
  assign _T_90629 = _T_90615[13]; // @[OneHot.scala 66:30:@39286.4]
  assign _T_90630 = _T_90615[14]; // @[OneHot.scala 66:30:@39287.4]
  assign _T_90631 = _T_90615[15]; // @[OneHot.scala 66:30:@39288.4]
  assign _T_90672 = loadRequest_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39306.4]
  assign _T_90673 = loadRequest_1 ? 16'h4000 : _T_90672; // @[Mux.scala 31:69:@39307.4]
  assign _T_90674 = loadRequest_0 ? 16'h2000 : _T_90673; // @[Mux.scala 31:69:@39308.4]
  assign _T_90675 = loadRequest_15 ? 16'h1000 : _T_90674; // @[Mux.scala 31:69:@39309.4]
  assign _T_90676 = loadRequest_14 ? 16'h800 : _T_90675; // @[Mux.scala 31:69:@39310.4]
  assign _T_90677 = loadRequest_13 ? 16'h400 : _T_90676; // @[Mux.scala 31:69:@39311.4]
  assign _T_90678 = loadRequest_12 ? 16'h200 : _T_90677; // @[Mux.scala 31:69:@39312.4]
  assign _T_90679 = loadRequest_11 ? 16'h100 : _T_90678; // @[Mux.scala 31:69:@39313.4]
  assign _T_90680 = loadRequest_10 ? 16'h80 : _T_90679; // @[Mux.scala 31:69:@39314.4]
  assign _T_90681 = loadRequest_9 ? 16'h40 : _T_90680; // @[Mux.scala 31:69:@39315.4]
  assign _T_90682 = loadRequest_8 ? 16'h20 : _T_90681; // @[Mux.scala 31:69:@39316.4]
  assign _T_90683 = loadRequest_7 ? 16'h10 : _T_90682; // @[Mux.scala 31:69:@39317.4]
  assign _T_90684 = loadRequest_6 ? 16'h8 : _T_90683; // @[Mux.scala 31:69:@39318.4]
  assign _T_90685 = loadRequest_5 ? 16'h4 : _T_90684; // @[Mux.scala 31:69:@39319.4]
  assign _T_90686 = loadRequest_4 ? 16'h2 : _T_90685; // @[Mux.scala 31:69:@39320.4]
  assign _T_90687 = loadRequest_3 ? 16'h1 : _T_90686; // @[Mux.scala 31:69:@39321.4]
  assign _T_90688 = _T_90687[0]; // @[OneHot.scala 66:30:@39322.4]
  assign _T_90689 = _T_90687[1]; // @[OneHot.scala 66:30:@39323.4]
  assign _T_90690 = _T_90687[2]; // @[OneHot.scala 66:30:@39324.4]
  assign _T_90691 = _T_90687[3]; // @[OneHot.scala 66:30:@39325.4]
  assign _T_90692 = _T_90687[4]; // @[OneHot.scala 66:30:@39326.4]
  assign _T_90693 = _T_90687[5]; // @[OneHot.scala 66:30:@39327.4]
  assign _T_90694 = _T_90687[6]; // @[OneHot.scala 66:30:@39328.4]
  assign _T_90695 = _T_90687[7]; // @[OneHot.scala 66:30:@39329.4]
  assign _T_90696 = _T_90687[8]; // @[OneHot.scala 66:30:@39330.4]
  assign _T_90697 = _T_90687[9]; // @[OneHot.scala 66:30:@39331.4]
  assign _T_90698 = _T_90687[10]; // @[OneHot.scala 66:30:@39332.4]
  assign _T_90699 = _T_90687[11]; // @[OneHot.scala 66:30:@39333.4]
  assign _T_90700 = _T_90687[12]; // @[OneHot.scala 66:30:@39334.4]
  assign _T_90701 = _T_90687[13]; // @[OneHot.scala 66:30:@39335.4]
  assign _T_90702 = _T_90687[14]; // @[OneHot.scala 66:30:@39336.4]
  assign _T_90703 = _T_90687[15]; // @[OneHot.scala 66:30:@39337.4]
  assign _T_90744 = loadRequest_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39355.4]
  assign _T_90745 = loadRequest_2 ? 16'h4000 : _T_90744; // @[Mux.scala 31:69:@39356.4]
  assign _T_90746 = loadRequest_1 ? 16'h2000 : _T_90745; // @[Mux.scala 31:69:@39357.4]
  assign _T_90747 = loadRequest_0 ? 16'h1000 : _T_90746; // @[Mux.scala 31:69:@39358.4]
  assign _T_90748 = loadRequest_15 ? 16'h800 : _T_90747; // @[Mux.scala 31:69:@39359.4]
  assign _T_90749 = loadRequest_14 ? 16'h400 : _T_90748; // @[Mux.scala 31:69:@39360.4]
  assign _T_90750 = loadRequest_13 ? 16'h200 : _T_90749; // @[Mux.scala 31:69:@39361.4]
  assign _T_90751 = loadRequest_12 ? 16'h100 : _T_90750; // @[Mux.scala 31:69:@39362.4]
  assign _T_90752 = loadRequest_11 ? 16'h80 : _T_90751; // @[Mux.scala 31:69:@39363.4]
  assign _T_90753 = loadRequest_10 ? 16'h40 : _T_90752; // @[Mux.scala 31:69:@39364.4]
  assign _T_90754 = loadRequest_9 ? 16'h20 : _T_90753; // @[Mux.scala 31:69:@39365.4]
  assign _T_90755 = loadRequest_8 ? 16'h10 : _T_90754; // @[Mux.scala 31:69:@39366.4]
  assign _T_90756 = loadRequest_7 ? 16'h8 : _T_90755; // @[Mux.scala 31:69:@39367.4]
  assign _T_90757 = loadRequest_6 ? 16'h4 : _T_90756; // @[Mux.scala 31:69:@39368.4]
  assign _T_90758 = loadRequest_5 ? 16'h2 : _T_90757; // @[Mux.scala 31:69:@39369.4]
  assign _T_90759 = loadRequest_4 ? 16'h1 : _T_90758; // @[Mux.scala 31:69:@39370.4]
  assign _T_90760 = _T_90759[0]; // @[OneHot.scala 66:30:@39371.4]
  assign _T_90761 = _T_90759[1]; // @[OneHot.scala 66:30:@39372.4]
  assign _T_90762 = _T_90759[2]; // @[OneHot.scala 66:30:@39373.4]
  assign _T_90763 = _T_90759[3]; // @[OneHot.scala 66:30:@39374.4]
  assign _T_90764 = _T_90759[4]; // @[OneHot.scala 66:30:@39375.4]
  assign _T_90765 = _T_90759[5]; // @[OneHot.scala 66:30:@39376.4]
  assign _T_90766 = _T_90759[6]; // @[OneHot.scala 66:30:@39377.4]
  assign _T_90767 = _T_90759[7]; // @[OneHot.scala 66:30:@39378.4]
  assign _T_90768 = _T_90759[8]; // @[OneHot.scala 66:30:@39379.4]
  assign _T_90769 = _T_90759[9]; // @[OneHot.scala 66:30:@39380.4]
  assign _T_90770 = _T_90759[10]; // @[OneHot.scala 66:30:@39381.4]
  assign _T_90771 = _T_90759[11]; // @[OneHot.scala 66:30:@39382.4]
  assign _T_90772 = _T_90759[12]; // @[OneHot.scala 66:30:@39383.4]
  assign _T_90773 = _T_90759[13]; // @[OneHot.scala 66:30:@39384.4]
  assign _T_90774 = _T_90759[14]; // @[OneHot.scala 66:30:@39385.4]
  assign _T_90775 = _T_90759[15]; // @[OneHot.scala 66:30:@39386.4]
  assign _T_90816 = loadRequest_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39404.4]
  assign _T_90817 = loadRequest_3 ? 16'h4000 : _T_90816; // @[Mux.scala 31:69:@39405.4]
  assign _T_90818 = loadRequest_2 ? 16'h2000 : _T_90817; // @[Mux.scala 31:69:@39406.4]
  assign _T_90819 = loadRequest_1 ? 16'h1000 : _T_90818; // @[Mux.scala 31:69:@39407.4]
  assign _T_90820 = loadRequest_0 ? 16'h800 : _T_90819; // @[Mux.scala 31:69:@39408.4]
  assign _T_90821 = loadRequest_15 ? 16'h400 : _T_90820; // @[Mux.scala 31:69:@39409.4]
  assign _T_90822 = loadRequest_14 ? 16'h200 : _T_90821; // @[Mux.scala 31:69:@39410.4]
  assign _T_90823 = loadRequest_13 ? 16'h100 : _T_90822; // @[Mux.scala 31:69:@39411.4]
  assign _T_90824 = loadRequest_12 ? 16'h80 : _T_90823; // @[Mux.scala 31:69:@39412.4]
  assign _T_90825 = loadRequest_11 ? 16'h40 : _T_90824; // @[Mux.scala 31:69:@39413.4]
  assign _T_90826 = loadRequest_10 ? 16'h20 : _T_90825; // @[Mux.scala 31:69:@39414.4]
  assign _T_90827 = loadRequest_9 ? 16'h10 : _T_90826; // @[Mux.scala 31:69:@39415.4]
  assign _T_90828 = loadRequest_8 ? 16'h8 : _T_90827; // @[Mux.scala 31:69:@39416.4]
  assign _T_90829 = loadRequest_7 ? 16'h4 : _T_90828; // @[Mux.scala 31:69:@39417.4]
  assign _T_90830 = loadRequest_6 ? 16'h2 : _T_90829; // @[Mux.scala 31:69:@39418.4]
  assign _T_90831 = loadRequest_5 ? 16'h1 : _T_90830; // @[Mux.scala 31:69:@39419.4]
  assign _T_90832 = _T_90831[0]; // @[OneHot.scala 66:30:@39420.4]
  assign _T_90833 = _T_90831[1]; // @[OneHot.scala 66:30:@39421.4]
  assign _T_90834 = _T_90831[2]; // @[OneHot.scala 66:30:@39422.4]
  assign _T_90835 = _T_90831[3]; // @[OneHot.scala 66:30:@39423.4]
  assign _T_90836 = _T_90831[4]; // @[OneHot.scala 66:30:@39424.4]
  assign _T_90837 = _T_90831[5]; // @[OneHot.scala 66:30:@39425.4]
  assign _T_90838 = _T_90831[6]; // @[OneHot.scala 66:30:@39426.4]
  assign _T_90839 = _T_90831[7]; // @[OneHot.scala 66:30:@39427.4]
  assign _T_90840 = _T_90831[8]; // @[OneHot.scala 66:30:@39428.4]
  assign _T_90841 = _T_90831[9]; // @[OneHot.scala 66:30:@39429.4]
  assign _T_90842 = _T_90831[10]; // @[OneHot.scala 66:30:@39430.4]
  assign _T_90843 = _T_90831[11]; // @[OneHot.scala 66:30:@39431.4]
  assign _T_90844 = _T_90831[12]; // @[OneHot.scala 66:30:@39432.4]
  assign _T_90845 = _T_90831[13]; // @[OneHot.scala 66:30:@39433.4]
  assign _T_90846 = _T_90831[14]; // @[OneHot.scala 66:30:@39434.4]
  assign _T_90847 = _T_90831[15]; // @[OneHot.scala 66:30:@39435.4]
  assign _T_90888 = loadRequest_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39453.4]
  assign _T_90889 = loadRequest_4 ? 16'h4000 : _T_90888; // @[Mux.scala 31:69:@39454.4]
  assign _T_90890 = loadRequest_3 ? 16'h2000 : _T_90889; // @[Mux.scala 31:69:@39455.4]
  assign _T_90891 = loadRequest_2 ? 16'h1000 : _T_90890; // @[Mux.scala 31:69:@39456.4]
  assign _T_90892 = loadRequest_1 ? 16'h800 : _T_90891; // @[Mux.scala 31:69:@39457.4]
  assign _T_90893 = loadRequest_0 ? 16'h400 : _T_90892; // @[Mux.scala 31:69:@39458.4]
  assign _T_90894 = loadRequest_15 ? 16'h200 : _T_90893; // @[Mux.scala 31:69:@39459.4]
  assign _T_90895 = loadRequest_14 ? 16'h100 : _T_90894; // @[Mux.scala 31:69:@39460.4]
  assign _T_90896 = loadRequest_13 ? 16'h80 : _T_90895; // @[Mux.scala 31:69:@39461.4]
  assign _T_90897 = loadRequest_12 ? 16'h40 : _T_90896; // @[Mux.scala 31:69:@39462.4]
  assign _T_90898 = loadRequest_11 ? 16'h20 : _T_90897; // @[Mux.scala 31:69:@39463.4]
  assign _T_90899 = loadRequest_10 ? 16'h10 : _T_90898; // @[Mux.scala 31:69:@39464.4]
  assign _T_90900 = loadRequest_9 ? 16'h8 : _T_90899; // @[Mux.scala 31:69:@39465.4]
  assign _T_90901 = loadRequest_8 ? 16'h4 : _T_90900; // @[Mux.scala 31:69:@39466.4]
  assign _T_90902 = loadRequest_7 ? 16'h2 : _T_90901; // @[Mux.scala 31:69:@39467.4]
  assign _T_90903 = loadRequest_6 ? 16'h1 : _T_90902; // @[Mux.scala 31:69:@39468.4]
  assign _T_90904 = _T_90903[0]; // @[OneHot.scala 66:30:@39469.4]
  assign _T_90905 = _T_90903[1]; // @[OneHot.scala 66:30:@39470.4]
  assign _T_90906 = _T_90903[2]; // @[OneHot.scala 66:30:@39471.4]
  assign _T_90907 = _T_90903[3]; // @[OneHot.scala 66:30:@39472.4]
  assign _T_90908 = _T_90903[4]; // @[OneHot.scala 66:30:@39473.4]
  assign _T_90909 = _T_90903[5]; // @[OneHot.scala 66:30:@39474.4]
  assign _T_90910 = _T_90903[6]; // @[OneHot.scala 66:30:@39475.4]
  assign _T_90911 = _T_90903[7]; // @[OneHot.scala 66:30:@39476.4]
  assign _T_90912 = _T_90903[8]; // @[OneHot.scala 66:30:@39477.4]
  assign _T_90913 = _T_90903[9]; // @[OneHot.scala 66:30:@39478.4]
  assign _T_90914 = _T_90903[10]; // @[OneHot.scala 66:30:@39479.4]
  assign _T_90915 = _T_90903[11]; // @[OneHot.scala 66:30:@39480.4]
  assign _T_90916 = _T_90903[12]; // @[OneHot.scala 66:30:@39481.4]
  assign _T_90917 = _T_90903[13]; // @[OneHot.scala 66:30:@39482.4]
  assign _T_90918 = _T_90903[14]; // @[OneHot.scala 66:30:@39483.4]
  assign _T_90919 = _T_90903[15]; // @[OneHot.scala 66:30:@39484.4]
  assign _T_90960 = loadRequest_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39502.4]
  assign _T_90961 = loadRequest_5 ? 16'h4000 : _T_90960; // @[Mux.scala 31:69:@39503.4]
  assign _T_90962 = loadRequest_4 ? 16'h2000 : _T_90961; // @[Mux.scala 31:69:@39504.4]
  assign _T_90963 = loadRequest_3 ? 16'h1000 : _T_90962; // @[Mux.scala 31:69:@39505.4]
  assign _T_90964 = loadRequest_2 ? 16'h800 : _T_90963; // @[Mux.scala 31:69:@39506.4]
  assign _T_90965 = loadRequest_1 ? 16'h400 : _T_90964; // @[Mux.scala 31:69:@39507.4]
  assign _T_90966 = loadRequest_0 ? 16'h200 : _T_90965; // @[Mux.scala 31:69:@39508.4]
  assign _T_90967 = loadRequest_15 ? 16'h100 : _T_90966; // @[Mux.scala 31:69:@39509.4]
  assign _T_90968 = loadRequest_14 ? 16'h80 : _T_90967; // @[Mux.scala 31:69:@39510.4]
  assign _T_90969 = loadRequest_13 ? 16'h40 : _T_90968; // @[Mux.scala 31:69:@39511.4]
  assign _T_90970 = loadRequest_12 ? 16'h20 : _T_90969; // @[Mux.scala 31:69:@39512.4]
  assign _T_90971 = loadRequest_11 ? 16'h10 : _T_90970; // @[Mux.scala 31:69:@39513.4]
  assign _T_90972 = loadRequest_10 ? 16'h8 : _T_90971; // @[Mux.scala 31:69:@39514.4]
  assign _T_90973 = loadRequest_9 ? 16'h4 : _T_90972; // @[Mux.scala 31:69:@39515.4]
  assign _T_90974 = loadRequest_8 ? 16'h2 : _T_90973; // @[Mux.scala 31:69:@39516.4]
  assign _T_90975 = loadRequest_7 ? 16'h1 : _T_90974; // @[Mux.scala 31:69:@39517.4]
  assign _T_90976 = _T_90975[0]; // @[OneHot.scala 66:30:@39518.4]
  assign _T_90977 = _T_90975[1]; // @[OneHot.scala 66:30:@39519.4]
  assign _T_90978 = _T_90975[2]; // @[OneHot.scala 66:30:@39520.4]
  assign _T_90979 = _T_90975[3]; // @[OneHot.scala 66:30:@39521.4]
  assign _T_90980 = _T_90975[4]; // @[OneHot.scala 66:30:@39522.4]
  assign _T_90981 = _T_90975[5]; // @[OneHot.scala 66:30:@39523.4]
  assign _T_90982 = _T_90975[6]; // @[OneHot.scala 66:30:@39524.4]
  assign _T_90983 = _T_90975[7]; // @[OneHot.scala 66:30:@39525.4]
  assign _T_90984 = _T_90975[8]; // @[OneHot.scala 66:30:@39526.4]
  assign _T_90985 = _T_90975[9]; // @[OneHot.scala 66:30:@39527.4]
  assign _T_90986 = _T_90975[10]; // @[OneHot.scala 66:30:@39528.4]
  assign _T_90987 = _T_90975[11]; // @[OneHot.scala 66:30:@39529.4]
  assign _T_90988 = _T_90975[12]; // @[OneHot.scala 66:30:@39530.4]
  assign _T_90989 = _T_90975[13]; // @[OneHot.scala 66:30:@39531.4]
  assign _T_90990 = _T_90975[14]; // @[OneHot.scala 66:30:@39532.4]
  assign _T_90991 = _T_90975[15]; // @[OneHot.scala 66:30:@39533.4]
  assign _T_91032 = loadRequest_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39551.4]
  assign _T_91033 = loadRequest_6 ? 16'h4000 : _T_91032; // @[Mux.scala 31:69:@39552.4]
  assign _T_91034 = loadRequest_5 ? 16'h2000 : _T_91033; // @[Mux.scala 31:69:@39553.4]
  assign _T_91035 = loadRequest_4 ? 16'h1000 : _T_91034; // @[Mux.scala 31:69:@39554.4]
  assign _T_91036 = loadRequest_3 ? 16'h800 : _T_91035; // @[Mux.scala 31:69:@39555.4]
  assign _T_91037 = loadRequest_2 ? 16'h400 : _T_91036; // @[Mux.scala 31:69:@39556.4]
  assign _T_91038 = loadRequest_1 ? 16'h200 : _T_91037; // @[Mux.scala 31:69:@39557.4]
  assign _T_91039 = loadRequest_0 ? 16'h100 : _T_91038; // @[Mux.scala 31:69:@39558.4]
  assign _T_91040 = loadRequest_15 ? 16'h80 : _T_91039; // @[Mux.scala 31:69:@39559.4]
  assign _T_91041 = loadRequest_14 ? 16'h40 : _T_91040; // @[Mux.scala 31:69:@39560.4]
  assign _T_91042 = loadRequest_13 ? 16'h20 : _T_91041; // @[Mux.scala 31:69:@39561.4]
  assign _T_91043 = loadRequest_12 ? 16'h10 : _T_91042; // @[Mux.scala 31:69:@39562.4]
  assign _T_91044 = loadRequest_11 ? 16'h8 : _T_91043; // @[Mux.scala 31:69:@39563.4]
  assign _T_91045 = loadRequest_10 ? 16'h4 : _T_91044; // @[Mux.scala 31:69:@39564.4]
  assign _T_91046 = loadRequest_9 ? 16'h2 : _T_91045; // @[Mux.scala 31:69:@39565.4]
  assign _T_91047 = loadRequest_8 ? 16'h1 : _T_91046; // @[Mux.scala 31:69:@39566.4]
  assign _T_91048 = _T_91047[0]; // @[OneHot.scala 66:30:@39567.4]
  assign _T_91049 = _T_91047[1]; // @[OneHot.scala 66:30:@39568.4]
  assign _T_91050 = _T_91047[2]; // @[OneHot.scala 66:30:@39569.4]
  assign _T_91051 = _T_91047[3]; // @[OneHot.scala 66:30:@39570.4]
  assign _T_91052 = _T_91047[4]; // @[OneHot.scala 66:30:@39571.4]
  assign _T_91053 = _T_91047[5]; // @[OneHot.scala 66:30:@39572.4]
  assign _T_91054 = _T_91047[6]; // @[OneHot.scala 66:30:@39573.4]
  assign _T_91055 = _T_91047[7]; // @[OneHot.scala 66:30:@39574.4]
  assign _T_91056 = _T_91047[8]; // @[OneHot.scala 66:30:@39575.4]
  assign _T_91057 = _T_91047[9]; // @[OneHot.scala 66:30:@39576.4]
  assign _T_91058 = _T_91047[10]; // @[OneHot.scala 66:30:@39577.4]
  assign _T_91059 = _T_91047[11]; // @[OneHot.scala 66:30:@39578.4]
  assign _T_91060 = _T_91047[12]; // @[OneHot.scala 66:30:@39579.4]
  assign _T_91061 = _T_91047[13]; // @[OneHot.scala 66:30:@39580.4]
  assign _T_91062 = _T_91047[14]; // @[OneHot.scala 66:30:@39581.4]
  assign _T_91063 = _T_91047[15]; // @[OneHot.scala 66:30:@39582.4]
  assign _T_91104 = loadRequest_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39600.4]
  assign _T_91105 = loadRequest_7 ? 16'h4000 : _T_91104; // @[Mux.scala 31:69:@39601.4]
  assign _T_91106 = loadRequest_6 ? 16'h2000 : _T_91105; // @[Mux.scala 31:69:@39602.4]
  assign _T_91107 = loadRequest_5 ? 16'h1000 : _T_91106; // @[Mux.scala 31:69:@39603.4]
  assign _T_91108 = loadRequest_4 ? 16'h800 : _T_91107; // @[Mux.scala 31:69:@39604.4]
  assign _T_91109 = loadRequest_3 ? 16'h400 : _T_91108; // @[Mux.scala 31:69:@39605.4]
  assign _T_91110 = loadRequest_2 ? 16'h200 : _T_91109; // @[Mux.scala 31:69:@39606.4]
  assign _T_91111 = loadRequest_1 ? 16'h100 : _T_91110; // @[Mux.scala 31:69:@39607.4]
  assign _T_91112 = loadRequest_0 ? 16'h80 : _T_91111; // @[Mux.scala 31:69:@39608.4]
  assign _T_91113 = loadRequest_15 ? 16'h40 : _T_91112; // @[Mux.scala 31:69:@39609.4]
  assign _T_91114 = loadRequest_14 ? 16'h20 : _T_91113; // @[Mux.scala 31:69:@39610.4]
  assign _T_91115 = loadRequest_13 ? 16'h10 : _T_91114; // @[Mux.scala 31:69:@39611.4]
  assign _T_91116 = loadRequest_12 ? 16'h8 : _T_91115; // @[Mux.scala 31:69:@39612.4]
  assign _T_91117 = loadRequest_11 ? 16'h4 : _T_91116; // @[Mux.scala 31:69:@39613.4]
  assign _T_91118 = loadRequest_10 ? 16'h2 : _T_91117; // @[Mux.scala 31:69:@39614.4]
  assign _T_91119 = loadRequest_9 ? 16'h1 : _T_91118; // @[Mux.scala 31:69:@39615.4]
  assign _T_91120 = _T_91119[0]; // @[OneHot.scala 66:30:@39616.4]
  assign _T_91121 = _T_91119[1]; // @[OneHot.scala 66:30:@39617.4]
  assign _T_91122 = _T_91119[2]; // @[OneHot.scala 66:30:@39618.4]
  assign _T_91123 = _T_91119[3]; // @[OneHot.scala 66:30:@39619.4]
  assign _T_91124 = _T_91119[4]; // @[OneHot.scala 66:30:@39620.4]
  assign _T_91125 = _T_91119[5]; // @[OneHot.scala 66:30:@39621.4]
  assign _T_91126 = _T_91119[6]; // @[OneHot.scala 66:30:@39622.4]
  assign _T_91127 = _T_91119[7]; // @[OneHot.scala 66:30:@39623.4]
  assign _T_91128 = _T_91119[8]; // @[OneHot.scala 66:30:@39624.4]
  assign _T_91129 = _T_91119[9]; // @[OneHot.scala 66:30:@39625.4]
  assign _T_91130 = _T_91119[10]; // @[OneHot.scala 66:30:@39626.4]
  assign _T_91131 = _T_91119[11]; // @[OneHot.scala 66:30:@39627.4]
  assign _T_91132 = _T_91119[12]; // @[OneHot.scala 66:30:@39628.4]
  assign _T_91133 = _T_91119[13]; // @[OneHot.scala 66:30:@39629.4]
  assign _T_91134 = _T_91119[14]; // @[OneHot.scala 66:30:@39630.4]
  assign _T_91135 = _T_91119[15]; // @[OneHot.scala 66:30:@39631.4]
  assign _T_91176 = loadRequest_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39649.4]
  assign _T_91177 = loadRequest_8 ? 16'h4000 : _T_91176; // @[Mux.scala 31:69:@39650.4]
  assign _T_91178 = loadRequest_7 ? 16'h2000 : _T_91177; // @[Mux.scala 31:69:@39651.4]
  assign _T_91179 = loadRequest_6 ? 16'h1000 : _T_91178; // @[Mux.scala 31:69:@39652.4]
  assign _T_91180 = loadRequest_5 ? 16'h800 : _T_91179; // @[Mux.scala 31:69:@39653.4]
  assign _T_91181 = loadRequest_4 ? 16'h400 : _T_91180; // @[Mux.scala 31:69:@39654.4]
  assign _T_91182 = loadRequest_3 ? 16'h200 : _T_91181; // @[Mux.scala 31:69:@39655.4]
  assign _T_91183 = loadRequest_2 ? 16'h100 : _T_91182; // @[Mux.scala 31:69:@39656.4]
  assign _T_91184 = loadRequest_1 ? 16'h80 : _T_91183; // @[Mux.scala 31:69:@39657.4]
  assign _T_91185 = loadRequest_0 ? 16'h40 : _T_91184; // @[Mux.scala 31:69:@39658.4]
  assign _T_91186 = loadRequest_15 ? 16'h20 : _T_91185; // @[Mux.scala 31:69:@39659.4]
  assign _T_91187 = loadRequest_14 ? 16'h10 : _T_91186; // @[Mux.scala 31:69:@39660.4]
  assign _T_91188 = loadRequest_13 ? 16'h8 : _T_91187; // @[Mux.scala 31:69:@39661.4]
  assign _T_91189 = loadRequest_12 ? 16'h4 : _T_91188; // @[Mux.scala 31:69:@39662.4]
  assign _T_91190 = loadRequest_11 ? 16'h2 : _T_91189; // @[Mux.scala 31:69:@39663.4]
  assign _T_91191 = loadRequest_10 ? 16'h1 : _T_91190; // @[Mux.scala 31:69:@39664.4]
  assign _T_91192 = _T_91191[0]; // @[OneHot.scala 66:30:@39665.4]
  assign _T_91193 = _T_91191[1]; // @[OneHot.scala 66:30:@39666.4]
  assign _T_91194 = _T_91191[2]; // @[OneHot.scala 66:30:@39667.4]
  assign _T_91195 = _T_91191[3]; // @[OneHot.scala 66:30:@39668.4]
  assign _T_91196 = _T_91191[4]; // @[OneHot.scala 66:30:@39669.4]
  assign _T_91197 = _T_91191[5]; // @[OneHot.scala 66:30:@39670.4]
  assign _T_91198 = _T_91191[6]; // @[OneHot.scala 66:30:@39671.4]
  assign _T_91199 = _T_91191[7]; // @[OneHot.scala 66:30:@39672.4]
  assign _T_91200 = _T_91191[8]; // @[OneHot.scala 66:30:@39673.4]
  assign _T_91201 = _T_91191[9]; // @[OneHot.scala 66:30:@39674.4]
  assign _T_91202 = _T_91191[10]; // @[OneHot.scala 66:30:@39675.4]
  assign _T_91203 = _T_91191[11]; // @[OneHot.scala 66:30:@39676.4]
  assign _T_91204 = _T_91191[12]; // @[OneHot.scala 66:30:@39677.4]
  assign _T_91205 = _T_91191[13]; // @[OneHot.scala 66:30:@39678.4]
  assign _T_91206 = _T_91191[14]; // @[OneHot.scala 66:30:@39679.4]
  assign _T_91207 = _T_91191[15]; // @[OneHot.scala 66:30:@39680.4]
  assign _T_91248 = loadRequest_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39698.4]
  assign _T_91249 = loadRequest_9 ? 16'h4000 : _T_91248; // @[Mux.scala 31:69:@39699.4]
  assign _T_91250 = loadRequest_8 ? 16'h2000 : _T_91249; // @[Mux.scala 31:69:@39700.4]
  assign _T_91251 = loadRequest_7 ? 16'h1000 : _T_91250; // @[Mux.scala 31:69:@39701.4]
  assign _T_91252 = loadRequest_6 ? 16'h800 : _T_91251; // @[Mux.scala 31:69:@39702.4]
  assign _T_91253 = loadRequest_5 ? 16'h400 : _T_91252; // @[Mux.scala 31:69:@39703.4]
  assign _T_91254 = loadRequest_4 ? 16'h200 : _T_91253; // @[Mux.scala 31:69:@39704.4]
  assign _T_91255 = loadRequest_3 ? 16'h100 : _T_91254; // @[Mux.scala 31:69:@39705.4]
  assign _T_91256 = loadRequest_2 ? 16'h80 : _T_91255; // @[Mux.scala 31:69:@39706.4]
  assign _T_91257 = loadRequest_1 ? 16'h40 : _T_91256; // @[Mux.scala 31:69:@39707.4]
  assign _T_91258 = loadRequest_0 ? 16'h20 : _T_91257; // @[Mux.scala 31:69:@39708.4]
  assign _T_91259 = loadRequest_15 ? 16'h10 : _T_91258; // @[Mux.scala 31:69:@39709.4]
  assign _T_91260 = loadRequest_14 ? 16'h8 : _T_91259; // @[Mux.scala 31:69:@39710.4]
  assign _T_91261 = loadRequest_13 ? 16'h4 : _T_91260; // @[Mux.scala 31:69:@39711.4]
  assign _T_91262 = loadRequest_12 ? 16'h2 : _T_91261; // @[Mux.scala 31:69:@39712.4]
  assign _T_91263 = loadRequest_11 ? 16'h1 : _T_91262; // @[Mux.scala 31:69:@39713.4]
  assign _T_91264 = _T_91263[0]; // @[OneHot.scala 66:30:@39714.4]
  assign _T_91265 = _T_91263[1]; // @[OneHot.scala 66:30:@39715.4]
  assign _T_91266 = _T_91263[2]; // @[OneHot.scala 66:30:@39716.4]
  assign _T_91267 = _T_91263[3]; // @[OneHot.scala 66:30:@39717.4]
  assign _T_91268 = _T_91263[4]; // @[OneHot.scala 66:30:@39718.4]
  assign _T_91269 = _T_91263[5]; // @[OneHot.scala 66:30:@39719.4]
  assign _T_91270 = _T_91263[6]; // @[OneHot.scala 66:30:@39720.4]
  assign _T_91271 = _T_91263[7]; // @[OneHot.scala 66:30:@39721.4]
  assign _T_91272 = _T_91263[8]; // @[OneHot.scala 66:30:@39722.4]
  assign _T_91273 = _T_91263[9]; // @[OneHot.scala 66:30:@39723.4]
  assign _T_91274 = _T_91263[10]; // @[OneHot.scala 66:30:@39724.4]
  assign _T_91275 = _T_91263[11]; // @[OneHot.scala 66:30:@39725.4]
  assign _T_91276 = _T_91263[12]; // @[OneHot.scala 66:30:@39726.4]
  assign _T_91277 = _T_91263[13]; // @[OneHot.scala 66:30:@39727.4]
  assign _T_91278 = _T_91263[14]; // @[OneHot.scala 66:30:@39728.4]
  assign _T_91279 = _T_91263[15]; // @[OneHot.scala 66:30:@39729.4]
  assign _T_91320 = loadRequest_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39747.4]
  assign _T_91321 = loadRequest_10 ? 16'h4000 : _T_91320; // @[Mux.scala 31:69:@39748.4]
  assign _T_91322 = loadRequest_9 ? 16'h2000 : _T_91321; // @[Mux.scala 31:69:@39749.4]
  assign _T_91323 = loadRequest_8 ? 16'h1000 : _T_91322; // @[Mux.scala 31:69:@39750.4]
  assign _T_91324 = loadRequest_7 ? 16'h800 : _T_91323; // @[Mux.scala 31:69:@39751.4]
  assign _T_91325 = loadRequest_6 ? 16'h400 : _T_91324; // @[Mux.scala 31:69:@39752.4]
  assign _T_91326 = loadRequest_5 ? 16'h200 : _T_91325; // @[Mux.scala 31:69:@39753.4]
  assign _T_91327 = loadRequest_4 ? 16'h100 : _T_91326; // @[Mux.scala 31:69:@39754.4]
  assign _T_91328 = loadRequest_3 ? 16'h80 : _T_91327; // @[Mux.scala 31:69:@39755.4]
  assign _T_91329 = loadRequest_2 ? 16'h40 : _T_91328; // @[Mux.scala 31:69:@39756.4]
  assign _T_91330 = loadRequest_1 ? 16'h20 : _T_91329; // @[Mux.scala 31:69:@39757.4]
  assign _T_91331 = loadRequest_0 ? 16'h10 : _T_91330; // @[Mux.scala 31:69:@39758.4]
  assign _T_91332 = loadRequest_15 ? 16'h8 : _T_91331; // @[Mux.scala 31:69:@39759.4]
  assign _T_91333 = loadRequest_14 ? 16'h4 : _T_91332; // @[Mux.scala 31:69:@39760.4]
  assign _T_91334 = loadRequest_13 ? 16'h2 : _T_91333; // @[Mux.scala 31:69:@39761.4]
  assign _T_91335 = loadRequest_12 ? 16'h1 : _T_91334; // @[Mux.scala 31:69:@39762.4]
  assign _T_91336 = _T_91335[0]; // @[OneHot.scala 66:30:@39763.4]
  assign _T_91337 = _T_91335[1]; // @[OneHot.scala 66:30:@39764.4]
  assign _T_91338 = _T_91335[2]; // @[OneHot.scala 66:30:@39765.4]
  assign _T_91339 = _T_91335[3]; // @[OneHot.scala 66:30:@39766.4]
  assign _T_91340 = _T_91335[4]; // @[OneHot.scala 66:30:@39767.4]
  assign _T_91341 = _T_91335[5]; // @[OneHot.scala 66:30:@39768.4]
  assign _T_91342 = _T_91335[6]; // @[OneHot.scala 66:30:@39769.4]
  assign _T_91343 = _T_91335[7]; // @[OneHot.scala 66:30:@39770.4]
  assign _T_91344 = _T_91335[8]; // @[OneHot.scala 66:30:@39771.4]
  assign _T_91345 = _T_91335[9]; // @[OneHot.scala 66:30:@39772.4]
  assign _T_91346 = _T_91335[10]; // @[OneHot.scala 66:30:@39773.4]
  assign _T_91347 = _T_91335[11]; // @[OneHot.scala 66:30:@39774.4]
  assign _T_91348 = _T_91335[12]; // @[OneHot.scala 66:30:@39775.4]
  assign _T_91349 = _T_91335[13]; // @[OneHot.scala 66:30:@39776.4]
  assign _T_91350 = _T_91335[14]; // @[OneHot.scala 66:30:@39777.4]
  assign _T_91351 = _T_91335[15]; // @[OneHot.scala 66:30:@39778.4]
  assign _T_91392 = loadRequest_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39796.4]
  assign _T_91393 = loadRequest_11 ? 16'h4000 : _T_91392; // @[Mux.scala 31:69:@39797.4]
  assign _T_91394 = loadRequest_10 ? 16'h2000 : _T_91393; // @[Mux.scala 31:69:@39798.4]
  assign _T_91395 = loadRequest_9 ? 16'h1000 : _T_91394; // @[Mux.scala 31:69:@39799.4]
  assign _T_91396 = loadRequest_8 ? 16'h800 : _T_91395; // @[Mux.scala 31:69:@39800.4]
  assign _T_91397 = loadRequest_7 ? 16'h400 : _T_91396; // @[Mux.scala 31:69:@39801.4]
  assign _T_91398 = loadRequest_6 ? 16'h200 : _T_91397; // @[Mux.scala 31:69:@39802.4]
  assign _T_91399 = loadRequest_5 ? 16'h100 : _T_91398; // @[Mux.scala 31:69:@39803.4]
  assign _T_91400 = loadRequest_4 ? 16'h80 : _T_91399; // @[Mux.scala 31:69:@39804.4]
  assign _T_91401 = loadRequest_3 ? 16'h40 : _T_91400; // @[Mux.scala 31:69:@39805.4]
  assign _T_91402 = loadRequest_2 ? 16'h20 : _T_91401; // @[Mux.scala 31:69:@39806.4]
  assign _T_91403 = loadRequest_1 ? 16'h10 : _T_91402; // @[Mux.scala 31:69:@39807.4]
  assign _T_91404 = loadRequest_0 ? 16'h8 : _T_91403; // @[Mux.scala 31:69:@39808.4]
  assign _T_91405 = loadRequest_15 ? 16'h4 : _T_91404; // @[Mux.scala 31:69:@39809.4]
  assign _T_91406 = loadRequest_14 ? 16'h2 : _T_91405; // @[Mux.scala 31:69:@39810.4]
  assign _T_91407 = loadRequest_13 ? 16'h1 : _T_91406; // @[Mux.scala 31:69:@39811.4]
  assign _T_91408 = _T_91407[0]; // @[OneHot.scala 66:30:@39812.4]
  assign _T_91409 = _T_91407[1]; // @[OneHot.scala 66:30:@39813.4]
  assign _T_91410 = _T_91407[2]; // @[OneHot.scala 66:30:@39814.4]
  assign _T_91411 = _T_91407[3]; // @[OneHot.scala 66:30:@39815.4]
  assign _T_91412 = _T_91407[4]; // @[OneHot.scala 66:30:@39816.4]
  assign _T_91413 = _T_91407[5]; // @[OneHot.scala 66:30:@39817.4]
  assign _T_91414 = _T_91407[6]; // @[OneHot.scala 66:30:@39818.4]
  assign _T_91415 = _T_91407[7]; // @[OneHot.scala 66:30:@39819.4]
  assign _T_91416 = _T_91407[8]; // @[OneHot.scala 66:30:@39820.4]
  assign _T_91417 = _T_91407[9]; // @[OneHot.scala 66:30:@39821.4]
  assign _T_91418 = _T_91407[10]; // @[OneHot.scala 66:30:@39822.4]
  assign _T_91419 = _T_91407[11]; // @[OneHot.scala 66:30:@39823.4]
  assign _T_91420 = _T_91407[12]; // @[OneHot.scala 66:30:@39824.4]
  assign _T_91421 = _T_91407[13]; // @[OneHot.scala 66:30:@39825.4]
  assign _T_91422 = _T_91407[14]; // @[OneHot.scala 66:30:@39826.4]
  assign _T_91423 = _T_91407[15]; // @[OneHot.scala 66:30:@39827.4]
  assign _T_91464 = loadRequest_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39845.4]
  assign _T_91465 = loadRequest_12 ? 16'h4000 : _T_91464; // @[Mux.scala 31:69:@39846.4]
  assign _T_91466 = loadRequest_11 ? 16'h2000 : _T_91465; // @[Mux.scala 31:69:@39847.4]
  assign _T_91467 = loadRequest_10 ? 16'h1000 : _T_91466; // @[Mux.scala 31:69:@39848.4]
  assign _T_91468 = loadRequest_9 ? 16'h800 : _T_91467; // @[Mux.scala 31:69:@39849.4]
  assign _T_91469 = loadRequest_8 ? 16'h400 : _T_91468; // @[Mux.scala 31:69:@39850.4]
  assign _T_91470 = loadRequest_7 ? 16'h200 : _T_91469; // @[Mux.scala 31:69:@39851.4]
  assign _T_91471 = loadRequest_6 ? 16'h100 : _T_91470; // @[Mux.scala 31:69:@39852.4]
  assign _T_91472 = loadRequest_5 ? 16'h80 : _T_91471; // @[Mux.scala 31:69:@39853.4]
  assign _T_91473 = loadRequest_4 ? 16'h40 : _T_91472; // @[Mux.scala 31:69:@39854.4]
  assign _T_91474 = loadRequest_3 ? 16'h20 : _T_91473; // @[Mux.scala 31:69:@39855.4]
  assign _T_91475 = loadRequest_2 ? 16'h10 : _T_91474; // @[Mux.scala 31:69:@39856.4]
  assign _T_91476 = loadRequest_1 ? 16'h8 : _T_91475; // @[Mux.scala 31:69:@39857.4]
  assign _T_91477 = loadRequest_0 ? 16'h4 : _T_91476; // @[Mux.scala 31:69:@39858.4]
  assign _T_91478 = loadRequest_15 ? 16'h2 : _T_91477; // @[Mux.scala 31:69:@39859.4]
  assign _T_91479 = loadRequest_14 ? 16'h1 : _T_91478; // @[Mux.scala 31:69:@39860.4]
  assign _T_91480 = _T_91479[0]; // @[OneHot.scala 66:30:@39861.4]
  assign _T_91481 = _T_91479[1]; // @[OneHot.scala 66:30:@39862.4]
  assign _T_91482 = _T_91479[2]; // @[OneHot.scala 66:30:@39863.4]
  assign _T_91483 = _T_91479[3]; // @[OneHot.scala 66:30:@39864.4]
  assign _T_91484 = _T_91479[4]; // @[OneHot.scala 66:30:@39865.4]
  assign _T_91485 = _T_91479[5]; // @[OneHot.scala 66:30:@39866.4]
  assign _T_91486 = _T_91479[6]; // @[OneHot.scala 66:30:@39867.4]
  assign _T_91487 = _T_91479[7]; // @[OneHot.scala 66:30:@39868.4]
  assign _T_91488 = _T_91479[8]; // @[OneHot.scala 66:30:@39869.4]
  assign _T_91489 = _T_91479[9]; // @[OneHot.scala 66:30:@39870.4]
  assign _T_91490 = _T_91479[10]; // @[OneHot.scala 66:30:@39871.4]
  assign _T_91491 = _T_91479[11]; // @[OneHot.scala 66:30:@39872.4]
  assign _T_91492 = _T_91479[12]; // @[OneHot.scala 66:30:@39873.4]
  assign _T_91493 = _T_91479[13]; // @[OneHot.scala 66:30:@39874.4]
  assign _T_91494 = _T_91479[14]; // @[OneHot.scala 66:30:@39875.4]
  assign _T_91495 = _T_91479[15]; // @[OneHot.scala 66:30:@39876.4]
  assign _T_91536 = loadRequest_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39894.4]
  assign _T_91537 = loadRequest_13 ? 16'h4000 : _T_91536; // @[Mux.scala 31:69:@39895.4]
  assign _T_91538 = loadRequest_12 ? 16'h2000 : _T_91537; // @[Mux.scala 31:69:@39896.4]
  assign _T_91539 = loadRequest_11 ? 16'h1000 : _T_91538; // @[Mux.scala 31:69:@39897.4]
  assign _T_91540 = loadRequest_10 ? 16'h800 : _T_91539; // @[Mux.scala 31:69:@39898.4]
  assign _T_91541 = loadRequest_9 ? 16'h400 : _T_91540; // @[Mux.scala 31:69:@39899.4]
  assign _T_91542 = loadRequest_8 ? 16'h200 : _T_91541; // @[Mux.scala 31:69:@39900.4]
  assign _T_91543 = loadRequest_7 ? 16'h100 : _T_91542; // @[Mux.scala 31:69:@39901.4]
  assign _T_91544 = loadRequest_6 ? 16'h80 : _T_91543; // @[Mux.scala 31:69:@39902.4]
  assign _T_91545 = loadRequest_5 ? 16'h40 : _T_91544; // @[Mux.scala 31:69:@39903.4]
  assign _T_91546 = loadRequest_4 ? 16'h20 : _T_91545; // @[Mux.scala 31:69:@39904.4]
  assign _T_91547 = loadRequest_3 ? 16'h10 : _T_91546; // @[Mux.scala 31:69:@39905.4]
  assign _T_91548 = loadRequest_2 ? 16'h8 : _T_91547; // @[Mux.scala 31:69:@39906.4]
  assign _T_91549 = loadRequest_1 ? 16'h4 : _T_91548; // @[Mux.scala 31:69:@39907.4]
  assign _T_91550 = loadRequest_0 ? 16'h2 : _T_91549; // @[Mux.scala 31:69:@39908.4]
  assign _T_91551 = loadRequest_15 ? 16'h1 : _T_91550; // @[Mux.scala 31:69:@39909.4]
  assign _T_91552 = _T_91551[0]; // @[OneHot.scala 66:30:@39910.4]
  assign _T_91553 = _T_91551[1]; // @[OneHot.scala 66:30:@39911.4]
  assign _T_91554 = _T_91551[2]; // @[OneHot.scala 66:30:@39912.4]
  assign _T_91555 = _T_91551[3]; // @[OneHot.scala 66:30:@39913.4]
  assign _T_91556 = _T_91551[4]; // @[OneHot.scala 66:30:@39914.4]
  assign _T_91557 = _T_91551[5]; // @[OneHot.scala 66:30:@39915.4]
  assign _T_91558 = _T_91551[6]; // @[OneHot.scala 66:30:@39916.4]
  assign _T_91559 = _T_91551[7]; // @[OneHot.scala 66:30:@39917.4]
  assign _T_91560 = _T_91551[8]; // @[OneHot.scala 66:30:@39918.4]
  assign _T_91561 = _T_91551[9]; // @[OneHot.scala 66:30:@39919.4]
  assign _T_91562 = _T_91551[10]; // @[OneHot.scala 66:30:@39920.4]
  assign _T_91563 = _T_91551[11]; // @[OneHot.scala 66:30:@39921.4]
  assign _T_91564 = _T_91551[12]; // @[OneHot.scala 66:30:@39922.4]
  assign _T_91565 = _T_91551[13]; // @[OneHot.scala 66:30:@39923.4]
  assign _T_91566 = _T_91551[14]; // @[OneHot.scala 66:30:@39924.4]
  assign _T_91567 = _T_91551[15]; // @[OneHot.scala 66:30:@39925.4]
  assign _T_91632 = {_T_90479,_T_90478,_T_90477,_T_90476,_T_90475,_T_90474,_T_90473,_T_90472}; // @[Mux.scala 19:72:@39949.4]
  assign _T_91640 = {_T_90487,_T_90486,_T_90485,_T_90484,_T_90483,_T_90482,_T_90481,_T_90480,_T_91632}; // @[Mux.scala 19:72:@39957.4]
  assign _T_91642 = _T_90400 ? _T_91640 : 16'h0; // @[Mux.scala 19:72:@39958.4]
  assign _T_91649 = {_T_90550,_T_90549,_T_90548,_T_90547,_T_90546,_T_90545,_T_90544,_T_90559}; // @[Mux.scala 19:72:@39965.4]
  assign _T_91657 = {_T_90558,_T_90557,_T_90556,_T_90555,_T_90554,_T_90553,_T_90552,_T_90551,_T_91649}; // @[Mux.scala 19:72:@39973.4]
  assign _T_91659 = _T_90401 ? _T_91657 : 16'h0; // @[Mux.scala 19:72:@39974.4]
  assign _T_91666 = {_T_90621,_T_90620,_T_90619,_T_90618,_T_90617,_T_90616,_T_90631,_T_90630}; // @[Mux.scala 19:72:@39981.4]
  assign _T_91674 = {_T_90629,_T_90628,_T_90627,_T_90626,_T_90625,_T_90624,_T_90623,_T_90622,_T_91666}; // @[Mux.scala 19:72:@39989.4]
  assign _T_91676 = _T_90402 ? _T_91674 : 16'h0; // @[Mux.scala 19:72:@39990.4]
  assign _T_91683 = {_T_90692,_T_90691,_T_90690,_T_90689,_T_90688,_T_90703,_T_90702,_T_90701}; // @[Mux.scala 19:72:@39997.4]
  assign _T_91691 = {_T_90700,_T_90699,_T_90698,_T_90697,_T_90696,_T_90695,_T_90694,_T_90693,_T_91683}; // @[Mux.scala 19:72:@40005.4]
  assign _T_91693 = _T_90403 ? _T_91691 : 16'h0; // @[Mux.scala 19:72:@40006.4]
  assign _T_91700 = {_T_90763,_T_90762,_T_90761,_T_90760,_T_90775,_T_90774,_T_90773,_T_90772}; // @[Mux.scala 19:72:@40013.4]
  assign _T_91708 = {_T_90771,_T_90770,_T_90769,_T_90768,_T_90767,_T_90766,_T_90765,_T_90764,_T_91700}; // @[Mux.scala 19:72:@40021.4]
  assign _T_91710 = _T_90404 ? _T_91708 : 16'h0; // @[Mux.scala 19:72:@40022.4]
  assign _T_91717 = {_T_90834,_T_90833,_T_90832,_T_90847,_T_90846,_T_90845,_T_90844,_T_90843}; // @[Mux.scala 19:72:@40029.4]
  assign _T_91725 = {_T_90842,_T_90841,_T_90840,_T_90839,_T_90838,_T_90837,_T_90836,_T_90835,_T_91717}; // @[Mux.scala 19:72:@40037.4]
  assign _T_91727 = _T_90405 ? _T_91725 : 16'h0; // @[Mux.scala 19:72:@40038.4]
  assign _T_91734 = {_T_90905,_T_90904,_T_90919,_T_90918,_T_90917,_T_90916,_T_90915,_T_90914}; // @[Mux.scala 19:72:@40045.4]
  assign _T_91742 = {_T_90913,_T_90912,_T_90911,_T_90910,_T_90909,_T_90908,_T_90907,_T_90906,_T_91734}; // @[Mux.scala 19:72:@40053.4]
  assign _T_91744 = _T_90406 ? _T_91742 : 16'h0; // @[Mux.scala 19:72:@40054.4]
  assign _T_91751 = {_T_90976,_T_90991,_T_90990,_T_90989,_T_90988,_T_90987,_T_90986,_T_90985}; // @[Mux.scala 19:72:@40061.4]
  assign _T_91759 = {_T_90984,_T_90983,_T_90982,_T_90981,_T_90980,_T_90979,_T_90978,_T_90977,_T_91751}; // @[Mux.scala 19:72:@40069.4]
  assign _T_91761 = _T_90407 ? _T_91759 : 16'h0; // @[Mux.scala 19:72:@40070.4]
  assign _T_91768 = {_T_91063,_T_91062,_T_91061,_T_91060,_T_91059,_T_91058,_T_91057,_T_91056}; // @[Mux.scala 19:72:@40077.4]
  assign _T_91776 = {_T_91055,_T_91054,_T_91053,_T_91052,_T_91051,_T_91050,_T_91049,_T_91048,_T_91768}; // @[Mux.scala 19:72:@40085.4]
  assign _T_91778 = _T_90408 ? _T_91776 : 16'h0; // @[Mux.scala 19:72:@40086.4]
  assign _T_91785 = {_T_91134,_T_91133,_T_91132,_T_91131,_T_91130,_T_91129,_T_91128,_T_91127}; // @[Mux.scala 19:72:@40093.4]
  assign _T_91793 = {_T_91126,_T_91125,_T_91124,_T_91123,_T_91122,_T_91121,_T_91120,_T_91135,_T_91785}; // @[Mux.scala 19:72:@40101.4]
  assign _T_91795 = _T_90409 ? _T_91793 : 16'h0; // @[Mux.scala 19:72:@40102.4]
  assign _T_91802 = {_T_91205,_T_91204,_T_91203,_T_91202,_T_91201,_T_91200,_T_91199,_T_91198}; // @[Mux.scala 19:72:@40109.4]
  assign _T_91810 = {_T_91197,_T_91196,_T_91195,_T_91194,_T_91193,_T_91192,_T_91207,_T_91206,_T_91802}; // @[Mux.scala 19:72:@40117.4]
  assign _T_91812 = _T_90410 ? _T_91810 : 16'h0; // @[Mux.scala 19:72:@40118.4]
  assign _T_91819 = {_T_91276,_T_91275,_T_91274,_T_91273,_T_91272,_T_91271,_T_91270,_T_91269}; // @[Mux.scala 19:72:@40125.4]
  assign _T_91827 = {_T_91268,_T_91267,_T_91266,_T_91265,_T_91264,_T_91279,_T_91278,_T_91277,_T_91819}; // @[Mux.scala 19:72:@40133.4]
  assign _T_91829 = _T_90411 ? _T_91827 : 16'h0; // @[Mux.scala 19:72:@40134.4]
  assign _T_91836 = {_T_91347,_T_91346,_T_91345,_T_91344,_T_91343,_T_91342,_T_91341,_T_91340}; // @[Mux.scala 19:72:@40141.4]
  assign _T_91844 = {_T_91339,_T_91338,_T_91337,_T_91336,_T_91351,_T_91350,_T_91349,_T_91348,_T_91836}; // @[Mux.scala 19:72:@40149.4]
  assign _T_91846 = _T_90412 ? _T_91844 : 16'h0; // @[Mux.scala 19:72:@40150.4]
  assign _T_91853 = {_T_91418,_T_91417,_T_91416,_T_91415,_T_91414,_T_91413,_T_91412,_T_91411}; // @[Mux.scala 19:72:@40157.4]
  assign _T_91861 = {_T_91410,_T_91409,_T_91408,_T_91423,_T_91422,_T_91421,_T_91420,_T_91419,_T_91853}; // @[Mux.scala 19:72:@40165.4]
  assign _T_91863 = _T_90413 ? _T_91861 : 16'h0; // @[Mux.scala 19:72:@40166.4]
  assign _T_91870 = {_T_91489,_T_91488,_T_91487,_T_91486,_T_91485,_T_91484,_T_91483,_T_91482}; // @[Mux.scala 19:72:@40173.4]
  assign _T_91878 = {_T_91481,_T_91480,_T_91495,_T_91494,_T_91493,_T_91492,_T_91491,_T_91490,_T_91870}; // @[Mux.scala 19:72:@40181.4]
  assign _T_91880 = _T_90414 ? _T_91878 : 16'h0; // @[Mux.scala 19:72:@40182.4]
  assign _T_91887 = {_T_91560,_T_91559,_T_91558,_T_91557,_T_91556,_T_91555,_T_91554,_T_91553}; // @[Mux.scala 19:72:@40189.4]
  assign _T_91895 = {_T_91552,_T_91567,_T_91566,_T_91565,_T_91564,_T_91563,_T_91562,_T_91561,_T_91887}; // @[Mux.scala 19:72:@40197.4]
  assign _T_91897 = _T_90415 ? _T_91895 : 16'h0; // @[Mux.scala 19:72:@40198.4]
  assign _T_91898 = _T_91642 | _T_91659; // @[Mux.scala 19:72:@40199.4]
  assign _T_91899 = _T_91898 | _T_91676; // @[Mux.scala 19:72:@40200.4]
  assign _T_91900 = _T_91899 | _T_91693; // @[Mux.scala 19:72:@40201.4]
  assign _T_91901 = _T_91900 | _T_91710; // @[Mux.scala 19:72:@40202.4]
  assign _T_91902 = _T_91901 | _T_91727; // @[Mux.scala 19:72:@40203.4]
  assign _T_91903 = _T_91902 | _T_91744; // @[Mux.scala 19:72:@40204.4]
  assign _T_91904 = _T_91903 | _T_91761; // @[Mux.scala 19:72:@40205.4]
  assign _T_91905 = _T_91904 | _T_91778; // @[Mux.scala 19:72:@40206.4]
  assign _T_91906 = _T_91905 | _T_91795; // @[Mux.scala 19:72:@40207.4]
  assign _T_91907 = _T_91906 | _T_91812; // @[Mux.scala 19:72:@40208.4]
  assign _T_91908 = _T_91907 | _T_91829; // @[Mux.scala 19:72:@40209.4]
  assign _T_91909 = _T_91908 | _T_91846; // @[Mux.scala 19:72:@40210.4]
  assign _T_91910 = _T_91909 | _T_91863; // @[Mux.scala 19:72:@40211.4]
  assign _T_91911 = _T_91910 | _T_91880; // @[Mux.scala 19:72:@40212.4]
  assign _T_91912 = _T_91911 | _T_91897; // @[Mux.scala 19:72:@40213.4]
  assign priorityLoadRequest_0 = _T_91912[0]; // @[Mux.scala 19:72:@40217.4]
  assign priorityLoadRequest_1 = _T_91912[1]; // @[Mux.scala 19:72:@40219.4]
  assign priorityLoadRequest_2 = _T_91912[2]; // @[Mux.scala 19:72:@40221.4]
  assign priorityLoadRequest_3 = _T_91912[3]; // @[Mux.scala 19:72:@40223.4]
  assign priorityLoadRequest_4 = _T_91912[4]; // @[Mux.scala 19:72:@40225.4]
  assign priorityLoadRequest_5 = _T_91912[5]; // @[Mux.scala 19:72:@40227.4]
  assign priorityLoadRequest_6 = _T_91912[6]; // @[Mux.scala 19:72:@40229.4]
  assign priorityLoadRequest_7 = _T_91912[7]; // @[Mux.scala 19:72:@40231.4]
  assign priorityLoadRequest_8 = _T_91912[8]; // @[Mux.scala 19:72:@40233.4]
  assign priorityLoadRequest_9 = _T_91912[9]; // @[Mux.scala 19:72:@40235.4]
  assign priorityLoadRequest_10 = _T_91912[10]; // @[Mux.scala 19:72:@40237.4]
  assign priorityLoadRequest_11 = _T_91912[11]; // @[Mux.scala 19:72:@40239.4]
  assign priorityLoadRequest_12 = _T_91912[12]; // @[Mux.scala 19:72:@40241.4]
  assign priorityLoadRequest_13 = _T_91912[13]; // @[Mux.scala 19:72:@40243.4]
  assign priorityLoadRequest_14 = _T_91912[14]; // @[Mux.scala 19:72:@40245.4]
  assign priorityLoadRequest_15 = _T_91912[15]; // @[Mux.scala 19:72:@40247.4]
  assign _GEN_1920 = io_memIsReadyForLoads ? priorityLoadRequest_0 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1921 = io_memIsReadyForLoads ? priorityLoadRequest_1 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1922 = io_memIsReadyForLoads ? priorityLoadRequest_2 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1923 = io_memIsReadyForLoads ? priorityLoadRequest_3 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1924 = io_memIsReadyForLoads ? priorityLoadRequest_4 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1925 = io_memIsReadyForLoads ? priorityLoadRequest_5 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1926 = io_memIsReadyForLoads ? priorityLoadRequest_6 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1927 = io_memIsReadyForLoads ? priorityLoadRequest_7 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1928 = io_memIsReadyForLoads ? priorityLoadRequest_8 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1929 = io_memIsReadyForLoads ? priorityLoadRequest_9 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1930 = io_memIsReadyForLoads ? priorityLoadRequest_10 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1931 = io_memIsReadyForLoads ? priorityLoadRequest_11 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1932 = io_memIsReadyForLoads ? priorityLoadRequest_12 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1933 = io_memIsReadyForLoads ? priorityLoadRequest_13 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1934 = io_memIsReadyForLoads ? priorityLoadRequest_14 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _GEN_1935 = io_memIsReadyForLoads ? priorityLoadRequest_15 : 1'h0; // @[LoadQueue.scala 208:31:@40267.4]
  assign _T_92307 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[LoadQueue.scala 238:58:@40485.8]
  assign _T_92315 = {storeAddrNotKnownFlagsPReg_0_15,storeAddrNotKnownFlagsPReg_0_14,storeAddrNotKnownFlagsPReg_0_13,storeAddrNotKnownFlagsPReg_0_12,storeAddrNotKnownFlagsPReg_0_11,storeAddrNotKnownFlagsPReg_0_10,storeAddrNotKnownFlagsPReg_0_9,storeAddrNotKnownFlagsPReg_0_8,_T_92307}; // @[LoadQueue.scala 238:58:@40493.8]
  assign _T_92322 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[LoadQueue.scala 238:96:@40500.8]
  assign _T_92330 = {lastConflict_0_15,lastConflict_0_14,lastConflict_0_13,lastConflict_0_12,lastConflict_0_11,lastConflict_0_10,lastConflict_0_9,lastConflict_0_8,_T_92322}; // @[LoadQueue.scala 238:96:@40508.8]
  assign _T_92331 = _T_92315 < _T_92330; // @[LoadQueue.scala 238:61:@40509.8]
  assign _T_92332 = canBypass_0 & _T_92331; // @[LoadQueue.scala 237:64:@40510.8]
  assign _GEN_1969 = _T_92261 ? _T_92332 : 1'h0; // @[LoadQueue.scala 230:110:@40442.6]
  assign bypassRequest_0 = _T_92253 ? _GEN_1969 : 1'h0; // @[LoadQueue.scala 229:71:@40436.4]
  assign _GEN_1936 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[LoadQueue.scala 217:34:@40324.6]
  assign _GEN_1937 = initBits_0 ? 1'h0 : _GEN_1936; // @[LoadQueue.scala 215:23:@40320.4]
  assign _T_92391 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[LoadQueue.scala 238:58:@40567.8]
  assign _T_92399 = {storeAddrNotKnownFlagsPReg_1_15,storeAddrNotKnownFlagsPReg_1_14,storeAddrNotKnownFlagsPReg_1_13,storeAddrNotKnownFlagsPReg_1_12,storeAddrNotKnownFlagsPReg_1_11,storeAddrNotKnownFlagsPReg_1_10,storeAddrNotKnownFlagsPReg_1_9,storeAddrNotKnownFlagsPReg_1_8,_T_92391}; // @[LoadQueue.scala 238:58:@40575.8]
  assign _T_92406 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[LoadQueue.scala 238:96:@40582.8]
  assign _T_92414 = {lastConflict_1_15,lastConflict_1_14,lastConflict_1_13,lastConflict_1_12,lastConflict_1_11,lastConflict_1_10,lastConflict_1_9,lastConflict_1_8,_T_92406}; // @[LoadQueue.scala 238:96:@40590.8]
  assign _T_92415 = _T_92399 < _T_92414; // @[LoadQueue.scala 238:61:@40591.8]
  assign _T_92416 = canBypass_1 & _T_92415; // @[LoadQueue.scala 237:64:@40592.8]
  assign _GEN_1973 = _T_92345 ? _T_92416 : 1'h0; // @[LoadQueue.scala 230:110:@40524.6]
  assign bypassRequest_1 = _T_92337 ? _GEN_1973 : 1'h0; // @[LoadQueue.scala 229:71:@40518.4]
  assign _GEN_1938 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[LoadQueue.scala 217:34:@40331.6]
  assign _GEN_1939 = initBits_1 ? 1'h0 : _GEN_1938; // @[LoadQueue.scala 215:23:@40327.4]
  assign _T_92475 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[LoadQueue.scala 238:58:@40649.8]
  assign _T_92483 = {storeAddrNotKnownFlagsPReg_2_15,storeAddrNotKnownFlagsPReg_2_14,storeAddrNotKnownFlagsPReg_2_13,storeAddrNotKnownFlagsPReg_2_12,storeAddrNotKnownFlagsPReg_2_11,storeAddrNotKnownFlagsPReg_2_10,storeAddrNotKnownFlagsPReg_2_9,storeAddrNotKnownFlagsPReg_2_8,_T_92475}; // @[LoadQueue.scala 238:58:@40657.8]
  assign _T_92490 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[LoadQueue.scala 238:96:@40664.8]
  assign _T_92498 = {lastConflict_2_15,lastConflict_2_14,lastConflict_2_13,lastConflict_2_12,lastConflict_2_11,lastConflict_2_10,lastConflict_2_9,lastConflict_2_8,_T_92490}; // @[LoadQueue.scala 238:96:@40672.8]
  assign _T_92499 = _T_92483 < _T_92498; // @[LoadQueue.scala 238:61:@40673.8]
  assign _T_92500 = canBypass_2 & _T_92499; // @[LoadQueue.scala 237:64:@40674.8]
  assign _GEN_1977 = _T_92429 ? _T_92500 : 1'h0; // @[LoadQueue.scala 230:110:@40606.6]
  assign bypassRequest_2 = _T_92421 ? _GEN_1977 : 1'h0; // @[LoadQueue.scala 229:71:@40600.4]
  assign _GEN_1940 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[LoadQueue.scala 217:34:@40338.6]
  assign _GEN_1941 = initBits_2 ? 1'h0 : _GEN_1940; // @[LoadQueue.scala 215:23:@40334.4]
  assign _T_92559 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[LoadQueue.scala 238:58:@40731.8]
  assign _T_92567 = {storeAddrNotKnownFlagsPReg_3_15,storeAddrNotKnownFlagsPReg_3_14,storeAddrNotKnownFlagsPReg_3_13,storeAddrNotKnownFlagsPReg_3_12,storeAddrNotKnownFlagsPReg_3_11,storeAddrNotKnownFlagsPReg_3_10,storeAddrNotKnownFlagsPReg_3_9,storeAddrNotKnownFlagsPReg_3_8,_T_92559}; // @[LoadQueue.scala 238:58:@40739.8]
  assign _T_92574 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[LoadQueue.scala 238:96:@40746.8]
  assign _T_92582 = {lastConflict_3_15,lastConflict_3_14,lastConflict_3_13,lastConflict_3_12,lastConflict_3_11,lastConflict_3_10,lastConflict_3_9,lastConflict_3_8,_T_92574}; // @[LoadQueue.scala 238:96:@40754.8]
  assign _T_92583 = _T_92567 < _T_92582; // @[LoadQueue.scala 238:61:@40755.8]
  assign _T_92584 = canBypass_3 & _T_92583; // @[LoadQueue.scala 237:64:@40756.8]
  assign _GEN_1981 = _T_92513 ? _T_92584 : 1'h0; // @[LoadQueue.scala 230:110:@40688.6]
  assign bypassRequest_3 = _T_92505 ? _GEN_1981 : 1'h0; // @[LoadQueue.scala 229:71:@40682.4]
  assign _GEN_1942 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[LoadQueue.scala 217:34:@40345.6]
  assign _GEN_1943 = initBits_3 ? 1'h0 : _GEN_1942; // @[LoadQueue.scala 215:23:@40341.4]
  assign _T_92643 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[LoadQueue.scala 238:58:@40813.8]
  assign _T_92651 = {storeAddrNotKnownFlagsPReg_4_15,storeAddrNotKnownFlagsPReg_4_14,storeAddrNotKnownFlagsPReg_4_13,storeAddrNotKnownFlagsPReg_4_12,storeAddrNotKnownFlagsPReg_4_11,storeAddrNotKnownFlagsPReg_4_10,storeAddrNotKnownFlagsPReg_4_9,storeAddrNotKnownFlagsPReg_4_8,_T_92643}; // @[LoadQueue.scala 238:58:@40821.8]
  assign _T_92658 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[LoadQueue.scala 238:96:@40828.8]
  assign _T_92666 = {lastConflict_4_15,lastConflict_4_14,lastConflict_4_13,lastConflict_4_12,lastConflict_4_11,lastConflict_4_10,lastConflict_4_9,lastConflict_4_8,_T_92658}; // @[LoadQueue.scala 238:96:@40836.8]
  assign _T_92667 = _T_92651 < _T_92666; // @[LoadQueue.scala 238:61:@40837.8]
  assign _T_92668 = canBypass_4 & _T_92667; // @[LoadQueue.scala 237:64:@40838.8]
  assign _GEN_1985 = _T_92597 ? _T_92668 : 1'h0; // @[LoadQueue.scala 230:110:@40770.6]
  assign bypassRequest_4 = _T_92589 ? _GEN_1985 : 1'h0; // @[LoadQueue.scala 229:71:@40764.4]
  assign _GEN_1944 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[LoadQueue.scala 217:34:@40352.6]
  assign _GEN_1945 = initBits_4 ? 1'h0 : _GEN_1944; // @[LoadQueue.scala 215:23:@40348.4]
  assign _T_92727 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[LoadQueue.scala 238:58:@40895.8]
  assign _T_92735 = {storeAddrNotKnownFlagsPReg_5_15,storeAddrNotKnownFlagsPReg_5_14,storeAddrNotKnownFlagsPReg_5_13,storeAddrNotKnownFlagsPReg_5_12,storeAddrNotKnownFlagsPReg_5_11,storeAddrNotKnownFlagsPReg_5_10,storeAddrNotKnownFlagsPReg_5_9,storeAddrNotKnownFlagsPReg_5_8,_T_92727}; // @[LoadQueue.scala 238:58:@40903.8]
  assign _T_92742 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[LoadQueue.scala 238:96:@40910.8]
  assign _T_92750 = {lastConflict_5_15,lastConflict_5_14,lastConflict_5_13,lastConflict_5_12,lastConflict_5_11,lastConflict_5_10,lastConflict_5_9,lastConflict_5_8,_T_92742}; // @[LoadQueue.scala 238:96:@40918.8]
  assign _T_92751 = _T_92735 < _T_92750; // @[LoadQueue.scala 238:61:@40919.8]
  assign _T_92752 = canBypass_5 & _T_92751; // @[LoadQueue.scala 237:64:@40920.8]
  assign _GEN_1989 = _T_92681 ? _T_92752 : 1'h0; // @[LoadQueue.scala 230:110:@40852.6]
  assign bypassRequest_5 = _T_92673 ? _GEN_1989 : 1'h0; // @[LoadQueue.scala 229:71:@40846.4]
  assign _GEN_1946 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[LoadQueue.scala 217:34:@40359.6]
  assign _GEN_1947 = initBits_5 ? 1'h0 : _GEN_1946; // @[LoadQueue.scala 215:23:@40355.4]
  assign _T_92811 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[LoadQueue.scala 238:58:@40977.8]
  assign _T_92819 = {storeAddrNotKnownFlagsPReg_6_15,storeAddrNotKnownFlagsPReg_6_14,storeAddrNotKnownFlagsPReg_6_13,storeAddrNotKnownFlagsPReg_6_12,storeAddrNotKnownFlagsPReg_6_11,storeAddrNotKnownFlagsPReg_6_10,storeAddrNotKnownFlagsPReg_6_9,storeAddrNotKnownFlagsPReg_6_8,_T_92811}; // @[LoadQueue.scala 238:58:@40985.8]
  assign _T_92826 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[LoadQueue.scala 238:96:@40992.8]
  assign _T_92834 = {lastConflict_6_15,lastConflict_6_14,lastConflict_6_13,lastConflict_6_12,lastConflict_6_11,lastConflict_6_10,lastConflict_6_9,lastConflict_6_8,_T_92826}; // @[LoadQueue.scala 238:96:@41000.8]
  assign _T_92835 = _T_92819 < _T_92834; // @[LoadQueue.scala 238:61:@41001.8]
  assign _T_92836 = canBypass_6 & _T_92835; // @[LoadQueue.scala 237:64:@41002.8]
  assign _GEN_1993 = _T_92765 ? _T_92836 : 1'h0; // @[LoadQueue.scala 230:110:@40934.6]
  assign bypassRequest_6 = _T_92757 ? _GEN_1993 : 1'h0; // @[LoadQueue.scala 229:71:@40928.4]
  assign _GEN_1948 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[LoadQueue.scala 217:34:@40366.6]
  assign _GEN_1949 = initBits_6 ? 1'h0 : _GEN_1948; // @[LoadQueue.scala 215:23:@40362.4]
  assign _T_92895 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[LoadQueue.scala 238:58:@41059.8]
  assign _T_92903 = {storeAddrNotKnownFlagsPReg_7_15,storeAddrNotKnownFlagsPReg_7_14,storeAddrNotKnownFlagsPReg_7_13,storeAddrNotKnownFlagsPReg_7_12,storeAddrNotKnownFlagsPReg_7_11,storeAddrNotKnownFlagsPReg_7_10,storeAddrNotKnownFlagsPReg_7_9,storeAddrNotKnownFlagsPReg_7_8,_T_92895}; // @[LoadQueue.scala 238:58:@41067.8]
  assign _T_92910 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[LoadQueue.scala 238:96:@41074.8]
  assign _T_92918 = {lastConflict_7_15,lastConflict_7_14,lastConflict_7_13,lastConflict_7_12,lastConflict_7_11,lastConflict_7_10,lastConflict_7_9,lastConflict_7_8,_T_92910}; // @[LoadQueue.scala 238:96:@41082.8]
  assign _T_92919 = _T_92903 < _T_92918; // @[LoadQueue.scala 238:61:@41083.8]
  assign _T_92920 = canBypass_7 & _T_92919; // @[LoadQueue.scala 237:64:@41084.8]
  assign _GEN_1997 = _T_92849 ? _T_92920 : 1'h0; // @[LoadQueue.scala 230:110:@41016.6]
  assign bypassRequest_7 = _T_92841 ? _GEN_1997 : 1'h0; // @[LoadQueue.scala 229:71:@41010.4]
  assign _GEN_1950 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[LoadQueue.scala 217:34:@40373.6]
  assign _GEN_1951 = initBits_7 ? 1'h0 : _GEN_1950; // @[LoadQueue.scala 215:23:@40369.4]
  assign _T_92979 = {storeAddrNotKnownFlagsPReg_8_7,storeAddrNotKnownFlagsPReg_8_6,storeAddrNotKnownFlagsPReg_8_5,storeAddrNotKnownFlagsPReg_8_4,storeAddrNotKnownFlagsPReg_8_3,storeAddrNotKnownFlagsPReg_8_2,storeAddrNotKnownFlagsPReg_8_1,storeAddrNotKnownFlagsPReg_8_0}; // @[LoadQueue.scala 238:58:@41141.8]
  assign _T_92987 = {storeAddrNotKnownFlagsPReg_8_15,storeAddrNotKnownFlagsPReg_8_14,storeAddrNotKnownFlagsPReg_8_13,storeAddrNotKnownFlagsPReg_8_12,storeAddrNotKnownFlagsPReg_8_11,storeAddrNotKnownFlagsPReg_8_10,storeAddrNotKnownFlagsPReg_8_9,storeAddrNotKnownFlagsPReg_8_8,_T_92979}; // @[LoadQueue.scala 238:58:@41149.8]
  assign _T_92994 = {lastConflict_8_7,lastConflict_8_6,lastConflict_8_5,lastConflict_8_4,lastConflict_8_3,lastConflict_8_2,lastConflict_8_1,lastConflict_8_0}; // @[LoadQueue.scala 238:96:@41156.8]
  assign _T_93002 = {lastConflict_8_15,lastConflict_8_14,lastConflict_8_13,lastConflict_8_12,lastConflict_8_11,lastConflict_8_10,lastConflict_8_9,lastConflict_8_8,_T_92994}; // @[LoadQueue.scala 238:96:@41164.8]
  assign _T_93003 = _T_92987 < _T_93002; // @[LoadQueue.scala 238:61:@41165.8]
  assign _T_93004 = canBypass_8 & _T_93003; // @[LoadQueue.scala 237:64:@41166.8]
  assign _GEN_2001 = _T_92933 ? _T_93004 : 1'h0; // @[LoadQueue.scala 230:110:@41098.6]
  assign bypassRequest_8 = _T_92925 ? _GEN_2001 : 1'h0; // @[LoadQueue.scala 229:71:@41092.4]
  assign _GEN_1952 = bypassRequest_8 ? 1'h1 : bypassInitiated_8; // @[LoadQueue.scala 217:34:@40380.6]
  assign _GEN_1953 = initBits_8 ? 1'h0 : _GEN_1952; // @[LoadQueue.scala 215:23:@40376.4]
  assign _T_93063 = {storeAddrNotKnownFlagsPReg_9_7,storeAddrNotKnownFlagsPReg_9_6,storeAddrNotKnownFlagsPReg_9_5,storeAddrNotKnownFlagsPReg_9_4,storeAddrNotKnownFlagsPReg_9_3,storeAddrNotKnownFlagsPReg_9_2,storeAddrNotKnownFlagsPReg_9_1,storeAddrNotKnownFlagsPReg_9_0}; // @[LoadQueue.scala 238:58:@41223.8]
  assign _T_93071 = {storeAddrNotKnownFlagsPReg_9_15,storeAddrNotKnownFlagsPReg_9_14,storeAddrNotKnownFlagsPReg_9_13,storeAddrNotKnownFlagsPReg_9_12,storeAddrNotKnownFlagsPReg_9_11,storeAddrNotKnownFlagsPReg_9_10,storeAddrNotKnownFlagsPReg_9_9,storeAddrNotKnownFlagsPReg_9_8,_T_93063}; // @[LoadQueue.scala 238:58:@41231.8]
  assign _T_93078 = {lastConflict_9_7,lastConflict_9_6,lastConflict_9_5,lastConflict_9_4,lastConflict_9_3,lastConflict_9_2,lastConflict_9_1,lastConflict_9_0}; // @[LoadQueue.scala 238:96:@41238.8]
  assign _T_93086 = {lastConflict_9_15,lastConflict_9_14,lastConflict_9_13,lastConflict_9_12,lastConflict_9_11,lastConflict_9_10,lastConflict_9_9,lastConflict_9_8,_T_93078}; // @[LoadQueue.scala 238:96:@41246.8]
  assign _T_93087 = _T_93071 < _T_93086; // @[LoadQueue.scala 238:61:@41247.8]
  assign _T_93088 = canBypass_9 & _T_93087; // @[LoadQueue.scala 237:64:@41248.8]
  assign _GEN_2005 = _T_93017 ? _T_93088 : 1'h0; // @[LoadQueue.scala 230:110:@41180.6]
  assign bypassRequest_9 = _T_93009 ? _GEN_2005 : 1'h0; // @[LoadQueue.scala 229:71:@41174.4]
  assign _GEN_1954 = bypassRequest_9 ? 1'h1 : bypassInitiated_9; // @[LoadQueue.scala 217:34:@40387.6]
  assign _GEN_1955 = initBits_9 ? 1'h0 : _GEN_1954; // @[LoadQueue.scala 215:23:@40383.4]
  assign _T_93147 = {storeAddrNotKnownFlagsPReg_10_7,storeAddrNotKnownFlagsPReg_10_6,storeAddrNotKnownFlagsPReg_10_5,storeAddrNotKnownFlagsPReg_10_4,storeAddrNotKnownFlagsPReg_10_3,storeAddrNotKnownFlagsPReg_10_2,storeAddrNotKnownFlagsPReg_10_1,storeAddrNotKnownFlagsPReg_10_0}; // @[LoadQueue.scala 238:58:@41305.8]
  assign _T_93155 = {storeAddrNotKnownFlagsPReg_10_15,storeAddrNotKnownFlagsPReg_10_14,storeAddrNotKnownFlagsPReg_10_13,storeAddrNotKnownFlagsPReg_10_12,storeAddrNotKnownFlagsPReg_10_11,storeAddrNotKnownFlagsPReg_10_10,storeAddrNotKnownFlagsPReg_10_9,storeAddrNotKnownFlagsPReg_10_8,_T_93147}; // @[LoadQueue.scala 238:58:@41313.8]
  assign _T_93162 = {lastConflict_10_7,lastConflict_10_6,lastConflict_10_5,lastConflict_10_4,lastConflict_10_3,lastConflict_10_2,lastConflict_10_1,lastConflict_10_0}; // @[LoadQueue.scala 238:96:@41320.8]
  assign _T_93170 = {lastConflict_10_15,lastConflict_10_14,lastConflict_10_13,lastConflict_10_12,lastConflict_10_11,lastConflict_10_10,lastConflict_10_9,lastConflict_10_8,_T_93162}; // @[LoadQueue.scala 238:96:@41328.8]
  assign _T_93171 = _T_93155 < _T_93170; // @[LoadQueue.scala 238:61:@41329.8]
  assign _T_93172 = canBypass_10 & _T_93171; // @[LoadQueue.scala 237:64:@41330.8]
  assign _GEN_2009 = _T_93101 ? _T_93172 : 1'h0; // @[LoadQueue.scala 230:110:@41262.6]
  assign bypassRequest_10 = _T_93093 ? _GEN_2009 : 1'h0; // @[LoadQueue.scala 229:71:@41256.4]
  assign _GEN_1956 = bypassRequest_10 ? 1'h1 : bypassInitiated_10; // @[LoadQueue.scala 217:34:@40394.6]
  assign _GEN_1957 = initBits_10 ? 1'h0 : _GEN_1956; // @[LoadQueue.scala 215:23:@40390.4]
  assign _T_93231 = {storeAddrNotKnownFlagsPReg_11_7,storeAddrNotKnownFlagsPReg_11_6,storeAddrNotKnownFlagsPReg_11_5,storeAddrNotKnownFlagsPReg_11_4,storeAddrNotKnownFlagsPReg_11_3,storeAddrNotKnownFlagsPReg_11_2,storeAddrNotKnownFlagsPReg_11_1,storeAddrNotKnownFlagsPReg_11_0}; // @[LoadQueue.scala 238:58:@41387.8]
  assign _T_93239 = {storeAddrNotKnownFlagsPReg_11_15,storeAddrNotKnownFlagsPReg_11_14,storeAddrNotKnownFlagsPReg_11_13,storeAddrNotKnownFlagsPReg_11_12,storeAddrNotKnownFlagsPReg_11_11,storeAddrNotKnownFlagsPReg_11_10,storeAddrNotKnownFlagsPReg_11_9,storeAddrNotKnownFlagsPReg_11_8,_T_93231}; // @[LoadQueue.scala 238:58:@41395.8]
  assign _T_93246 = {lastConflict_11_7,lastConflict_11_6,lastConflict_11_5,lastConflict_11_4,lastConflict_11_3,lastConflict_11_2,lastConflict_11_1,lastConflict_11_0}; // @[LoadQueue.scala 238:96:@41402.8]
  assign _T_93254 = {lastConflict_11_15,lastConflict_11_14,lastConflict_11_13,lastConflict_11_12,lastConflict_11_11,lastConflict_11_10,lastConflict_11_9,lastConflict_11_8,_T_93246}; // @[LoadQueue.scala 238:96:@41410.8]
  assign _T_93255 = _T_93239 < _T_93254; // @[LoadQueue.scala 238:61:@41411.8]
  assign _T_93256 = canBypass_11 & _T_93255; // @[LoadQueue.scala 237:64:@41412.8]
  assign _GEN_2013 = _T_93185 ? _T_93256 : 1'h0; // @[LoadQueue.scala 230:110:@41344.6]
  assign bypassRequest_11 = _T_93177 ? _GEN_2013 : 1'h0; // @[LoadQueue.scala 229:71:@41338.4]
  assign _GEN_1958 = bypassRequest_11 ? 1'h1 : bypassInitiated_11; // @[LoadQueue.scala 217:34:@40401.6]
  assign _GEN_1959 = initBits_11 ? 1'h0 : _GEN_1958; // @[LoadQueue.scala 215:23:@40397.4]
  assign _T_93315 = {storeAddrNotKnownFlagsPReg_12_7,storeAddrNotKnownFlagsPReg_12_6,storeAddrNotKnownFlagsPReg_12_5,storeAddrNotKnownFlagsPReg_12_4,storeAddrNotKnownFlagsPReg_12_3,storeAddrNotKnownFlagsPReg_12_2,storeAddrNotKnownFlagsPReg_12_1,storeAddrNotKnownFlagsPReg_12_0}; // @[LoadQueue.scala 238:58:@41469.8]
  assign _T_93323 = {storeAddrNotKnownFlagsPReg_12_15,storeAddrNotKnownFlagsPReg_12_14,storeAddrNotKnownFlagsPReg_12_13,storeAddrNotKnownFlagsPReg_12_12,storeAddrNotKnownFlagsPReg_12_11,storeAddrNotKnownFlagsPReg_12_10,storeAddrNotKnownFlagsPReg_12_9,storeAddrNotKnownFlagsPReg_12_8,_T_93315}; // @[LoadQueue.scala 238:58:@41477.8]
  assign _T_93330 = {lastConflict_12_7,lastConflict_12_6,lastConflict_12_5,lastConflict_12_4,lastConflict_12_3,lastConflict_12_2,lastConflict_12_1,lastConflict_12_0}; // @[LoadQueue.scala 238:96:@41484.8]
  assign _T_93338 = {lastConflict_12_15,lastConflict_12_14,lastConflict_12_13,lastConflict_12_12,lastConflict_12_11,lastConflict_12_10,lastConflict_12_9,lastConflict_12_8,_T_93330}; // @[LoadQueue.scala 238:96:@41492.8]
  assign _T_93339 = _T_93323 < _T_93338; // @[LoadQueue.scala 238:61:@41493.8]
  assign _T_93340 = canBypass_12 & _T_93339; // @[LoadQueue.scala 237:64:@41494.8]
  assign _GEN_2017 = _T_93269 ? _T_93340 : 1'h0; // @[LoadQueue.scala 230:110:@41426.6]
  assign bypassRequest_12 = _T_93261 ? _GEN_2017 : 1'h0; // @[LoadQueue.scala 229:71:@41420.4]
  assign _GEN_1960 = bypassRequest_12 ? 1'h1 : bypassInitiated_12; // @[LoadQueue.scala 217:34:@40408.6]
  assign _GEN_1961 = initBits_12 ? 1'h0 : _GEN_1960; // @[LoadQueue.scala 215:23:@40404.4]
  assign _T_93399 = {storeAddrNotKnownFlagsPReg_13_7,storeAddrNotKnownFlagsPReg_13_6,storeAddrNotKnownFlagsPReg_13_5,storeAddrNotKnownFlagsPReg_13_4,storeAddrNotKnownFlagsPReg_13_3,storeAddrNotKnownFlagsPReg_13_2,storeAddrNotKnownFlagsPReg_13_1,storeAddrNotKnownFlagsPReg_13_0}; // @[LoadQueue.scala 238:58:@41551.8]
  assign _T_93407 = {storeAddrNotKnownFlagsPReg_13_15,storeAddrNotKnownFlagsPReg_13_14,storeAddrNotKnownFlagsPReg_13_13,storeAddrNotKnownFlagsPReg_13_12,storeAddrNotKnownFlagsPReg_13_11,storeAddrNotKnownFlagsPReg_13_10,storeAddrNotKnownFlagsPReg_13_9,storeAddrNotKnownFlagsPReg_13_8,_T_93399}; // @[LoadQueue.scala 238:58:@41559.8]
  assign _T_93414 = {lastConflict_13_7,lastConflict_13_6,lastConflict_13_5,lastConflict_13_4,lastConflict_13_3,lastConflict_13_2,lastConflict_13_1,lastConflict_13_0}; // @[LoadQueue.scala 238:96:@41566.8]
  assign _T_93422 = {lastConflict_13_15,lastConflict_13_14,lastConflict_13_13,lastConflict_13_12,lastConflict_13_11,lastConflict_13_10,lastConflict_13_9,lastConflict_13_8,_T_93414}; // @[LoadQueue.scala 238:96:@41574.8]
  assign _T_93423 = _T_93407 < _T_93422; // @[LoadQueue.scala 238:61:@41575.8]
  assign _T_93424 = canBypass_13 & _T_93423; // @[LoadQueue.scala 237:64:@41576.8]
  assign _GEN_2021 = _T_93353 ? _T_93424 : 1'h0; // @[LoadQueue.scala 230:110:@41508.6]
  assign bypassRequest_13 = _T_93345 ? _GEN_2021 : 1'h0; // @[LoadQueue.scala 229:71:@41502.4]
  assign _GEN_1962 = bypassRequest_13 ? 1'h1 : bypassInitiated_13; // @[LoadQueue.scala 217:34:@40415.6]
  assign _GEN_1963 = initBits_13 ? 1'h0 : _GEN_1962; // @[LoadQueue.scala 215:23:@40411.4]
  assign _T_93483 = {storeAddrNotKnownFlagsPReg_14_7,storeAddrNotKnownFlagsPReg_14_6,storeAddrNotKnownFlagsPReg_14_5,storeAddrNotKnownFlagsPReg_14_4,storeAddrNotKnownFlagsPReg_14_3,storeAddrNotKnownFlagsPReg_14_2,storeAddrNotKnownFlagsPReg_14_1,storeAddrNotKnownFlagsPReg_14_0}; // @[LoadQueue.scala 238:58:@41633.8]
  assign _T_93491 = {storeAddrNotKnownFlagsPReg_14_15,storeAddrNotKnownFlagsPReg_14_14,storeAddrNotKnownFlagsPReg_14_13,storeAddrNotKnownFlagsPReg_14_12,storeAddrNotKnownFlagsPReg_14_11,storeAddrNotKnownFlagsPReg_14_10,storeAddrNotKnownFlagsPReg_14_9,storeAddrNotKnownFlagsPReg_14_8,_T_93483}; // @[LoadQueue.scala 238:58:@41641.8]
  assign _T_93498 = {lastConflict_14_7,lastConflict_14_6,lastConflict_14_5,lastConflict_14_4,lastConflict_14_3,lastConflict_14_2,lastConflict_14_1,lastConflict_14_0}; // @[LoadQueue.scala 238:96:@41648.8]
  assign _T_93506 = {lastConflict_14_15,lastConflict_14_14,lastConflict_14_13,lastConflict_14_12,lastConflict_14_11,lastConflict_14_10,lastConflict_14_9,lastConflict_14_8,_T_93498}; // @[LoadQueue.scala 238:96:@41656.8]
  assign _T_93507 = _T_93491 < _T_93506; // @[LoadQueue.scala 238:61:@41657.8]
  assign _T_93508 = canBypass_14 & _T_93507; // @[LoadQueue.scala 237:64:@41658.8]
  assign _GEN_2025 = _T_93437 ? _T_93508 : 1'h0; // @[LoadQueue.scala 230:110:@41590.6]
  assign bypassRequest_14 = _T_93429 ? _GEN_2025 : 1'h0; // @[LoadQueue.scala 229:71:@41584.4]
  assign _GEN_1964 = bypassRequest_14 ? 1'h1 : bypassInitiated_14; // @[LoadQueue.scala 217:34:@40422.6]
  assign _GEN_1965 = initBits_14 ? 1'h0 : _GEN_1964; // @[LoadQueue.scala 215:23:@40418.4]
  assign _T_93567 = {storeAddrNotKnownFlagsPReg_15_7,storeAddrNotKnownFlagsPReg_15_6,storeAddrNotKnownFlagsPReg_15_5,storeAddrNotKnownFlagsPReg_15_4,storeAddrNotKnownFlagsPReg_15_3,storeAddrNotKnownFlagsPReg_15_2,storeAddrNotKnownFlagsPReg_15_1,storeAddrNotKnownFlagsPReg_15_0}; // @[LoadQueue.scala 238:58:@41715.8]
  assign _T_93575 = {storeAddrNotKnownFlagsPReg_15_15,storeAddrNotKnownFlagsPReg_15_14,storeAddrNotKnownFlagsPReg_15_13,storeAddrNotKnownFlagsPReg_15_12,storeAddrNotKnownFlagsPReg_15_11,storeAddrNotKnownFlagsPReg_15_10,storeAddrNotKnownFlagsPReg_15_9,storeAddrNotKnownFlagsPReg_15_8,_T_93567}; // @[LoadQueue.scala 238:58:@41723.8]
  assign _T_93582 = {lastConflict_15_7,lastConflict_15_6,lastConflict_15_5,lastConflict_15_4,lastConflict_15_3,lastConflict_15_2,lastConflict_15_1,lastConflict_15_0}; // @[LoadQueue.scala 238:96:@41730.8]
  assign _T_93590 = {lastConflict_15_15,lastConflict_15_14,lastConflict_15_13,lastConflict_15_12,lastConflict_15_11,lastConflict_15_10,lastConflict_15_9,lastConflict_15_8,_T_93582}; // @[LoadQueue.scala 238:96:@41738.8]
  assign _T_93591 = _T_93575 < _T_93590; // @[LoadQueue.scala 238:61:@41739.8]
  assign _T_93592 = canBypass_15 & _T_93591; // @[LoadQueue.scala 237:64:@41740.8]
  assign _GEN_2029 = _T_93521 ? _T_93592 : 1'h0; // @[LoadQueue.scala 230:110:@41672.6]
  assign bypassRequest_15 = _T_93513 ? _GEN_2029 : 1'h0; // @[LoadQueue.scala 229:71:@41666.4]
  assign _GEN_1966 = bypassRequest_15 ? 1'h1 : bypassInitiated_15; // @[LoadQueue.scala 217:34:@40429.6]
  assign _GEN_1967 = initBits_15 ? 1'h0 : _GEN_1966; // @[LoadQueue.scala 215:23:@40425.4]
  assign _T_93596 = loadRequest_0 | loadRequest_1; // @[LoadQueue.scala 247:28:@41746.4]
  assign _T_93597 = _T_93596 | loadRequest_2; // @[LoadQueue.scala 247:28:@41747.4]
  assign _T_93598 = _T_93597 | loadRequest_3; // @[LoadQueue.scala 247:28:@41748.4]
  assign _T_93599 = _T_93598 | loadRequest_4; // @[LoadQueue.scala 247:28:@41749.4]
  assign _T_93600 = _T_93599 | loadRequest_5; // @[LoadQueue.scala 247:28:@41750.4]
  assign _T_93601 = _T_93600 | loadRequest_6; // @[LoadQueue.scala 247:28:@41751.4]
  assign _T_93602 = _T_93601 | loadRequest_7; // @[LoadQueue.scala 247:28:@41752.4]
  assign _T_93603 = _T_93602 | loadRequest_8; // @[LoadQueue.scala 247:28:@41753.4]
  assign _T_93604 = _T_93603 | loadRequest_9; // @[LoadQueue.scala 247:28:@41754.4]
  assign _T_93605 = _T_93604 | loadRequest_10; // @[LoadQueue.scala 247:28:@41755.4]
  assign _T_93606 = _T_93605 | loadRequest_11; // @[LoadQueue.scala 247:28:@41756.4]
  assign _T_93607 = _T_93606 | loadRequest_12; // @[LoadQueue.scala 247:28:@41757.4]
  assign _T_93608 = _T_93607 | loadRequest_13; // @[LoadQueue.scala 247:28:@41758.4]
  assign _T_93609 = _T_93608 | loadRequest_14; // @[LoadQueue.scala 247:28:@41759.4]
  assign _T_93610 = _T_93609 | loadRequest_15; // @[LoadQueue.scala 247:28:@41760.4]
  assign _T_93627 = priorityLoadRequest_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@41762.6]
  assign _T_93628 = priorityLoadRequest_13 ? 4'hd : _T_93627; // @[Mux.scala 31:69:@41763.6]
  assign _T_93629 = priorityLoadRequest_12 ? 4'hc : _T_93628; // @[Mux.scala 31:69:@41764.6]
  assign _T_93630 = priorityLoadRequest_11 ? 4'hb : _T_93629; // @[Mux.scala 31:69:@41765.6]
  assign _T_93631 = priorityLoadRequest_10 ? 4'ha : _T_93630; // @[Mux.scala 31:69:@41766.6]
  assign _T_93632 = priorityLoadRequest_9 ? 4'h9 : _T_93631; // @[Mux.scala 31:69:@41767.6]
  assign _T_93633 = priorityLoadRequest_8 ? 4'h8 : _T_93632; // @[Mux.scala 31:69:@41768.6]
  assign _T_93634 = priorityLoadRequest_7 ? 4'h7 : _T_93633; // @[Mux.scala 31:69:@41769.6]
  assign _T_93635 = priorityLoadRequest_6 ? 4'h6 : _T_93634; // @[Mux.scala 31:69:@41770.6]
  assign _T_93636 = priorityLoadRequest_5 ? 4'h5 : _T_93635; // @[Mux.scala 31:69:@41771.6]
  assign _T_93637 = priorityLoadRequest_4 ? 4'h4 : _T_93636; // @[Mux.scala 31:69:@41772.6]
  assign _T_93638 = priorityLoadRequest_3 ? 4'h3 : _T_93637; // @[Mux.scala 31:69:@41773.6]
  assign _T_93639 = priorityLoadRequest_2 ? 4'h2 : _T_93638; // @[Mux.scala 31:69:@41774.6]
  assign _T_93640 = priorityLoadRequest_1 ? 4'h1 : _T_93639; // @[Mux.scala 31:69:@41775.6]
  assign _T_93641 = priorityLoadRequest_0 ? 4'h0 : _T_93640; // @[Mux.scala 31:69:@41776.6]
  assign _GEN_2033 = 4'h1 == _T_93641 ? addrQ_1 : addrQ_0; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2034 = 4'h2 == _T_93641 ? addrQ_2 : _GEN_2033; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2035 = 4'h3 == _T_93641 ? addrQ_3 : _GEN_2034; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2036 = 4'h4 == _T_93641 ? addrQ_4 : _GEN_2035; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2037 = 4'h5 == _T_93641 ? addrQ_5 : _GEN_2036; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2038 = 4'h6 == _T_93641 ? addrQ_6 : _GEN_2037; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2039 = 4'h7 == _T_93641 ? addrQ_7 : _GEN_2038; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2040 = 4'h8 == _T_93641 ? addrQ_8 : _GEN_2039; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2041 = 4'h9 == _T_93641 ? addrQ_9 : _GEN_2040; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2042 = 4'ha == _T_93641 ? addrQ_10 : _GEN_2041; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2043 = 4'hb == _T_93641 ? addrQ_11 : _GEN_2042; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2044 = 4'hc == _T_93641 ? addrQ_12 : _GEN_2043; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2045 = 4'hd == _T_93641 ? addrQ_13 : _GEN_2044; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2046 = 4'he == _T_93641 ? addrQ_14 : _GEN_2045; // @[LoadQueue.scala 248:24:@41777.6]
  assign _GEN_2047 = 4'hf == _T_93641 ? addrQ_15 : _GEN_2046; // @[LoadQueue.scala 248:24:@41777.6]
  assign _T_93649 = prevPriorityRequest_0 | bypassRequest_0; // @[LoadQueue.scala 261:41:@41788.6]
  assign _GEN_2050 = _T_93649 ? 1'h1 : dataKnown_0; // @[LoadQueue.scala 261:62:@41789.6]
  assign _GEN_2051 = initBits_0 ? 1'h0 : _GEN_2050; // @[LoadQueue.scala 259:25:@41784.4]
  assign _T_93652 = prevPriorityRequest_1 | bypassRequest_1; // @[LoadQueue.scala 261:41:@41796.6]
  assign _GEN_2052 = _T_93652 ? 1'h1 : dataKnown_1; // @[LoadQueue.scala 261:62:@41797.6]
  assign _GEN_2053 = initBits_1 ? 1'h0 : _GEN_2052; // @[LoadQueue.scala 259:25:@41792.4]
  assign _T_93655 = prevPriorityRequest_2 | bypassRequest_2; // @[LoadQueue.scala 261:41:@41804.6]
  assign _GEN_2054 = _T_93655 ? 1'h1 : dataKnown_2; // @[LoadQueue.scala 261:62:@41805.6]
  assign _GEN_2055 = initBits_2 ? 1'h0 : _GEN_2054; // @[LoadQueue.scala 259:25:@41800.4]
  assign _T_93658 = prevPriorityRequest_3 | bypassRequest_3; // @[LoadQueue.scala 261:41:@41812.6]
  assign _GEN_2056 = _T_93658 ? 1'h1 : dataKnown_3; // @[LoadQueue.scala 261:62:@41813.6]
  assign _GEN_2057 = initBits_3 ? 1'h0 : _GEN_2056; // @[LoadQueue.scala 259:25:@41808.4]
  assign _T_93661 = prevPriorityRequest_4 | bypassRequest_4; // @[LoadQueue.scala 261:41:@41820.6]
  assign _GEN_2058 = _T_93661 ? 1'h1 : dataKnown_4; // @[LoadQueue.scala 261:62:@41821.6]
  assign _GEN_2059 = initBits_4 ? 1'h0 : _GEN_2058; // @[LoadQueue.scala 259:25:@41816.4]
  assign _T_93664 = prevPriorityRequest_5 | bypassRequest_5; // @[LoadQueue.scala 261:41:@41828.6]
  assign _GEN_2060 = _T_93664 ? 1'h1 : dataKnown_5; // @[LoadQueue.scala 261:62:@41829.6]
  assign _GEN_2061 = initBits_5 ? 1'h0 : _GEN_2060; // @[LoadQueue.scala 259:25:@41824.4]
  assign _T_93667 = prevPriorityRequest_6 | bypassRequest_6; // @[LoadQueue.scala 261:41:@41836.6]
  assign _GEN_2062 = _T_93667 ? 1'h1 : dataKnown_6; // @[LoadQueue.scala 261:62:@41837.6]
  assign _GEN_2063 = initBits_6 ? 1'h0 : _GEN_2062; // @[LoadQueue.scala 259:25:@41832.4]
  assign _T_93670 = prevPriorityRequest_7 | bypassRequest_7; // @[LoadQueue.scala 261:41:@41844.6]
  assign _GEN_2064 = _T_93670 ? 1'h1 : dataKnown_7; // @[LoadQueue.scala 261:62:@41845.6]
  assign _GEN_2065 = initBits_7 ? 1'h0 : _GEN_2064; // @[LoadQueue.scala 259:25:@41840.4]
  assign _T_93673 = prevPriorityRequest_8 | bypassRequest_8; // @[LoadQueue.scala 261:41:@41852.6]
  assign _GEN_2066 = _T_93673 ? 1'h1 : dataKnown_8; // @[LoadQueue.scala 261:62:@41853.6]
  assign _GEN_2067 = initBits_8 ? 1'h0 : _GEN_2066; // @[LoadQueue.scala 259:25:@41848.4]
  assign _T_93676 = prevPriorityRequest_9 | bypassRequest_9; // @[LoadQueue.scala 261:41:@41860.6]
  assign _GEN_2068 = _T_93676 ? 1'h1 : dataKnown_9; // @[LoadQueue.scala 261:62:@41861.6]
  assign _GEN_2069 = initBits_9 ? 1'h0 : _GEN_2068; // @[LoadQueue.scala 259:25:@41856.4]
  assign _T_93679 = prevPriorityRequest_10 | bypassRequest_10; // @[LoadQueue.scala 261:41:@41868.6]
  assign _GEN_2070 = _T_93679 ? 1'h1 : dataKnown_10; // @[LoadQueue.scala 261:62:@41869.6]
  assign _GEN_2071 = initBits_10 ? 1'h0 : _GEN_2070; // @[LoadQueue.scala 259:25:@41864.4]
  assign _T_93682 = prevPriorityRequest_11 | bypassRequest_11; // @[LoadQueue.scala 261:41:@41876.6]
  assign _GEN_2072 = _T_93682 ? 1'h1 : dataKnown_11; // @[LoadQueue.scala 261:62:@41877.6]
  assign _GEN_2073 = initBits_11 ? 1'h0 : _GEN_2072; // @[LoadQueue.scala 259:25:@41872.4]
  assign _T_93685 = prevPriorityRequest_12 | bypassRequest_12; // @[LoadQueue.scala 261:41:@41884.6]
  assign _GEN_2074 = _T_93685 ? 1'h1 : dataKnown_12; // @[LoadQueue.scala 261:62:@41885.6]
  assign _GEN_2075 = initBits_12 ? 1'h0 : _GEN_2074; // @[LoadQueue.scala 259:25:@41880.4]
  assign _T_93688 = prevPriorityRequest_13 | bypassRequest_13; // @[LoadQueue.scala 261:41:@41892.6]
  assign _GEN_2076 = _T_93688 ? 1'h1 : dataKnown_13; // @[LoadQueue.scala 261:62:@41893.6]
  assign _GEN_2077 = initBits_13 ? 1'h0 : _GEN_2076; // @[LoadQueue.scala 259:25:@41888.4]
  assign _T_93691 = prevPriorityRequest_14 | bypassRequest_14; // @[LoadQueue.scala 261:41:@41900.6]
  assign _GEN_2078 = _T_93691 ? 1'h1 : dataKnown_14; // @[LoadQueue.scala 261:62:@41901.6]
  assign _GEN_2079 = initBits_14 ? 1'h0 : _GEN_2078; // @[LoadQueue.scala 259:25:@41896.4]
  assign _T_93694 = prevPriorityRequest_15 | bypassRequest_15; // @[LoadQueue.scala 261:41:@41908.6]
  assign _GEN_2080 = _T_93694 ? 1'h1 : dataKnown_15; // @[LoadQueue.scala 261:62:@41909.6]
  assign _GEN_2081 = initBits_15 ? 1'h0 : _GEN_2080; // @[LoadQueue.scala 259:25:@41904.4]
  assign _GEN_2082 = prevPriorityRequest_0 ? io_loadDataFromMem : dataQ_0; // @[LoadQueue.scala 269:44:@41916.6]
  assign _GEN_2083 = bypassRequest_0 ? bypassVal_0 : _GEN_2082; // @[LoadQueue.scala 267:32:@41912.4]
  assign _GEN_2084 = prevPriorityRequest_1 ? io_loadDataFromMem : dataQ_1; // @[LoadQueue.scala 269:44:@41923.6]
  assign _GEN_2085 = bypassRequest_1 ? bypassVal_1 : _GEN_2084; // @[LoadQueue.scala 267:32:@41919.4]
  assign _GEN_2086 = prevPriorityRequest_2 ? io_loadDataFromMem : dataQ_2; // @[LoadQueue.scala 269:44:@41930.6]
  assign _GEN_2087 = bypassRequest_2 ? bypassVal_2 : _GEN_2086; // @[LoadQueue.scala 267:32:@41926.4]
  assign _GEN_2088 = prevPriorityRequest_3 ? io_loadDataFromMem : dataQ_3; // @[LoadQueue.scala 269:44:@41937.6]
  assign _GEN_2089 = bypassRequest_3 ? bypassVal_3 : _GEN_2088; // @[LoadQueue.scala 267:32:@41933.4]
  assign _GEN_2090 = prevPriorityRequest_4 ? io_loadDataFromMem : dataQ_4; // @[LoadQueue.scala 269:44:@41944.6]
  assign _GEN_2091 = bypassRequest_4 ? bypassVal_4 : _GEN_2090; // @[LoadQueue.scala 267:32:@41940.4]
  assign _GEN_2092 = prevPriorityRequest_5 ? io_loadDataFromMem : dataQ_5; // @[LoadQueue.scala 269:44:@41951.6]
  assign _GEN_2093 = bypassRequest_5 ? bypassVal_5 : _GEN_2092; // @[LoadQueue.scala 267:32:@41947.4]
  assign _GEN_2094 = prevPriorityRequest_6 ? io_loadDataFromMem : dataQ_6; // @[LoadQueue.scala 269:44:@41958.6]
  assign _GEN_2095 = bypassRequest_6 ? bypassVal_6 : _GEN_2094; // @[LoadQueue.scala 267:32:@41954.4]
  assign _GEN_2096 = prevPriorityRequest_7 ? io_loadDataFromMem : dataQ_7; // @[LoadQueue.scala 269:44:@41965.6]
  assign _GEN_2097 = bypassRequest_7 ? bypassVal_7 : _GEN_2096; // @[LoadQueue.scala 267:32:@41961.4]
  assign _GEN_2098 = prevPriorityRequest_8 ? io_loadDataFromMem : dataQ_8; // @[LoadQueue.scala 269:44:@41972.6]
  assign _GEN_2099 = bypassRequest_8 ? bypassVal_8 : _GEN_2098; // @[LoadQueue.scala 267:32:@41968.4]
  assign _GEN_2100 = prevPriorityRequest_9 ? io_loadDataFromMem : dataQ_9; // @[LoadQueue.scala 269:44:@41979.6]
  assign _GEN_2101 = bypassRequest_9 ? bypassVal_9 : _GEN_2100; // @[LoadQueue.scala 267:32:@41975.4]
  assign _GEN_2102 = prevPriorityRequest_10 ? io_loadDataFromMem : dataQ_10; // @[LoadQueue.scala 269:44:@41986.6]
  assign _GEN_2103 = bypassRequest_10 ? bypassVal_10 : _GEN_2102; // @[LoadQueue.scala 267:32:@41982.4]
  assign _GEN_2104 = prevPriorityRequest_11 ? io_loadDataFromMem : dataQ_11; // @[LoadQueue.scala 269:44:@41993.6]
  assign _GEN_2105 = bypassRequest_11 ? bypassVal_11 : _GEN_2104; // @[LoadQueue.scala 267:32:@41989.4]
  assign _GEN_2106 = prevPriorityRequest_12 ? io_loadDataFromMem : dataQ_12; // @[LoadQueue.scala 269:44:@42000.6]
  assign _GEN_2107 = bypassRequest_12 ? bypassVal_12 : _GEN_2106; // @[LoadQueue.scala 267:32:@41996.4]
  assign _GEN_2108 = prevPriorityRequest_13 ? io_loadDataFromMem : dataQ_13; // @[LoadQueue.scala 269:44:@42007.6]
  assign _GEN_2109 = bypassRequest_13 ? bypassVal_13 : _GEN_2108; // @[LoadQueue.scala 267:32:@42003.4]
  assign _GEN_2110 = prevPriorityRequest_14 ? io_loadDataFromMem : dataQ_14; // @[LoadQueue.scala 269:44:@42014.6]
  assign _GEN_2111 = bypassRequest_14 ? bypassVal_14 : _GEN_2110; // @[LoadQueue.scala 267:32:@42010.4]
  assign _GEN_2112 = prevPriorityRequest_15 ? io_loadDataFromMem : dataQ_15; // @[LoadQueue.scala 269:44:@42021.6]
  assign _GEN_2113 = bypassRequest_15 ? bypassVal_15 : _GEN_2112; // @[LoadQueue.scala 267:32:@42017.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[LoadQueue.scala 286:69:@42025.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[LoadQueue.scala 286:69:@42027.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[LoadQueue.scala 286:69:@42029.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[LoadQueue.scala 286:69:@42031.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[LoadQueue.scala 286:69:@42033.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[LoadQueue.scala 286:69:@42035.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[LoadQueue.scala 286:69:@42037.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[LoadQueue.scala 286:69:@42039.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[LoadQueue.scala 286:69:@42041.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[LoadQueue.scala 286:69:@42043.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[LoadQueue.scala 286:69:@42045.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[LoadQueue.scala 286:69:@42047.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[LoadQueue.scala 286:69:@42049.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[LoadQueue.scala 286:69:@42051.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[LoadQueue.scala 286:69:@42053.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[LoadQueue.scala 286:69:@42055.4]
  assign _T_94179 = addrKnown_0 == 1'h0; // @[LoadQueue.scala 298:86:@42059.4]
  assign _T_94180 = entriesPorts_0_0 & _T_94179; // @[LoadQueue.scala 298:83:@42060.4]
  assign _T_94182 = addrKnown_1 == 1'h0; // @[LoadQueue.scala 298:86:@42061.4]
  assign _T_94183 = entriesPorts_0_1 & _T_94182; // @[LoadQueue.scala 298:83:@42062.4]
  assign _T_94185 = addrKnown_2 == 1'h0; // @[LoadQueue.scala 298:86:@42063.4]
  assign _T_94186 = entriesPorts_0_2 & _T_94185; // @[LoadQueue.scala 298:83:@42064.4]
  assign _T_94188 = addrKnown_3 == 1'h0; // @[LoadQueue.scala 298:86:@42065.4]
  assign _T_94189 = entriesPorts_0_3 & _T_94188; // @[LoadQueue.scala 298:83:@42066.4]
  assign _T_94191 = addrKnown_4 == 1'h0; // @[LoadQueue.scala 298:86:@42067.4]
  assign _T_94192 = entriesPorts_0_4 & _T_94191; // @[LoadQueue.scala 298:83:@42068.4]
  assign _T_94194 = addrKnown_5 == 1'h0; // @[LoadQueue.scala 298:86:@42069.4]
  assign _T_94195 = entriesPorts_0_5 & _T_94194; // @[LoadQueue.scala 298:83:@42070.4]
  assign _T_94197 = addrKnown_6 == 1'h0; // @[LoadQueue.scala 298:86:@42071.4]
  assign _T_94198 = entriesPorts_0_6 & _T_94197; // @[LoadQueue.scala 298:83:@42072.4]
  assign _T_94200 = addrKnown_7 == 1'h0; // @[LoadQueue.scala 298:86:@42073.4]
  assign _T_94201 = entriesPorts_0_7 & _T_94200; // @[LoadQueue.scala 298:83:@42074.4]
  assign _T_94203 = addrKnown_8 == 1'h0; // @[LoadQueue.scala 298:86:@42075.4]
  assign _T_94204 = entriesPorts_0_8 & _T_94203; // @[LoadQueue.scala 298:83:@42076.4]
  assign _T_94206 = addrKnown_9 == 1'h0; // @[LoadQueue.scala 298:86:@42077.4]
  assign _T_94207 = entriesPorts_0_9 & _T_94206; // @[LoadQueue.scala 298:83:@42078.4]
  assign _T_94209 = addrKnown_10 == 1'h0; // @[LoadQueue.scala 298:86:@42079.4]
  assign _T_94210 = entriesPorts_0_10 & _T_94209; // @[LoadQueue.scala 298:83:@42080.4]
  assign _T_94212 = addrKnown_11 == 1'h0; // @[LoadQueue.scala 298:86:@42081.4]
  assign _T_94213 = entriesPorts_0_11 & _T_94212; // @[LoadQueue.scala 298:83:@42082.4]
  assign _T_94215 = addrKnown_12 == 1'h0; // @[LoadQueue.scala 298:86:@42083.4]
  assign _T_94216 = entriesPorts_0_12 & _T_94215; // @[LoadQueue.scala 298:83:@42084.4]
  assign _T_94218 = addrKnown_13 == 1'h0; // @[LoadQueue.scala 298:86:@42085.4]
  assign _T_94219 = entriesPorts_0_13 & _T_94218; // @[LoadQueue.scala 298:83:@42086.4]
  assign _T_94221 = addrKnown_14 == 1'h0; // @[LoadQueue.scala 298:86:@42087.4]
  assign _T_94222 = entriesPorts_0_14 & _T_94221; // @[LoadQueue.scala 298:83:@42088.4]
  assign _T_94224 = addrKnown_15 == 1'h0; // @[LoadQueue.scala 298:86:@42089.4]
  assign _T_94225 = entriesPorts_0_15 & _T_94224; // @[LoadQueue.scala 298:83:@42090.4]
  assign _T_94308 = _T_94225 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42144.4]
  assign _T_94309 = _T_94222 ? 16'h4000 : _T_94308; // @[Mux.scala 31:69:@42145.4]
  assign _T_94310 = _T_94219 ? 16'h2000 : _T_94309; // @[Mux.scala 31:69:@42146.4]
  assign _T_94311 = _T_94216 ? 16'h1000 : _T_94310; // @[Mux.scala 31:69:@42147.4]
  assign _T_94312 = _T_94213 ? 16'h800 : _T_94311; // @[Mux.scala 31:69:@42148.4]
  assign _T_94313 = _T_94210 ? 16'h400 : _T_94312; // @[Mux.scala 31:69:@42149.4]
  assign _T_94314 = _T_94207 ? 16'h200 : _T_94313; // @[Mux.scala 31:69:@42150.4]
  assign _T_94315 = _T_94204 ? 16'h100 : _T_94314; // @[Mux.scala 31:69:@42151.4]
  assign _T_94316 = _T_94201 ? 16'h80 : _T_94315; // @[Mux.scala 31:69:@42152.4]
  assign _T_94317 = _T_94198 ? 16'h40 : _T_94316; // @[Mux.scala 31:69:@42153.4]
  assign _T_94318 = _T_94195 ? 16'h20 : _T_94317; // @[Mux.scala 31:69:@42154.4]
  assign _T_94319 = _T_94192 ? 16'h10 : _T_94318; // @[Mux.scala 31:69:@42155.4]
  assign _T_94320 = _T_94189 ? 16'h8 : _T_94319; // @[Mux.scala 31:69:@42156.4]
  assign _T_94321 = _T_94186 ? 16'h4 : _T_94320; // @[Mux.scala 31:69:@42157.4]
  assign _T_94322 = _T_94183 ? 16'h2 : _T_94321; // @[Mux.scala 31:69:@42158.4]
  assign _T_94323 = _T_94180 ? 16'h1 : _T_94322; // @[Mux.scala 31:69:@42159.4]
  assign _T_94324 = _T_94323[0]; // @[OneHot.scala 66:30:@42160.4]
  assign _T_94325 = _T_94323[1]; // @[OneHot.scala 66:30:@42161.4]
  assign _T_94326 = _T_94323[2]; // @[OneHot.scala 66:30:@42162.4]
  assign _T_94327 = _T_94323[3]; // @[OneHot.scala 66:30:@42163.4]
  assign _T_94328 = _T_94323[4]; // @[OneHot.scala 66:30:@42164.4]
  assign _T_94329 = _T_94323[5]; // @[OneHot.scala 66:30:@42165.4]
  assign _T_94330 = _T_94323[6]; // @[OneHot.scala 66:30:@42166.4]
  assign _T_94331 = _T_94323[7]; // @[OneHot.scala 66:30:@42167.4]
  assign _T_94332 = _T_94323[8]; // @[OneHot.scala 66:30:@42168.4]
  assign _T_94333 = _T_94323[9]; // @[OneHot.scala 66:30:@42169.4]
  assign _T_94334 = _T_94323[10]; // @[OneHot.scala 66:30:@42170.4]
  assign _T_94335 = _T_94323[11]; // @[OneHot.scala 66:30:@42171.4]
  assign _T_94336 = _T_94323[12]; // @[OneHot.scala 66:30:@42172.4]
  assign _T_94337 = _T_94323[13]; // @[OneHot.scala 66:30:@42173.4]
  assign _T_94338 = _T_94323[14]; // @[OneHot.scala 66:30:@42174.4]
  assign _T_94339 = _T_94323[15]; // @[OneHot.scala 66:30:@42175.4]
  assign _T_94380 = _T_94180 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42193.4]
  assign _T_94381 = _T_94225 ? 16'h4000 : _T_94380; // @[Mux.scala 31:69:@42194.4]
  assign _T_94382 = _T_94222 ? 16'h2000 : _T_94381; // @[Mux.scala 31:69:@42195.4]
  assign _T_94383 = _T_94219 ? 16'h1000 : _T_94382; // @[Mux.scala 31:69:@42196.4]
  assign _T_94384 = _T_94216 ? 16'h800 : _T_94383; // @[Mux.scala 31:69:@42197.4]
  assign _T_94385 = _T_94213 ? 16'h400 : _T_94384; // @[Mux.scala 31:69:@42198.4]
  assign _T_94386 = _T_94210 ? 16'h200 : _T_94385; // @[Mux.scala 31:69:@42199.4]
  assign _T_94387 = _T_94207 ? 16'h100 : _T_94386; // @[Mux.scala 31:69:@42200.4]
  assign _T_94388 = _T_94204 ? 16'h80 : _T_94387; // @[Mux.scala 31:69:@42201.4]
  assign _T_94389 = _T_94201 ? 16'h40 : _T_94388; // @[Mux.scala 31:69:@42202.4]
  assign _T_94390 = _T_94198 ? 16'h20 : _T_94389; // @[Mux.scala 31:69:@42203.4]
  assign _T_94391 = _T_94195 ? 16'h10 : _T_94390; // @[Mux.scala 31:69:@42204.4]
  assign _T_94392 = _T_94192 ? 16'h8 : _T_94391; // @[Mux.scala 31:69:@42205.4]
  assign _T_94393 = _T_94189 ? 16'h4 : _T_94392; // @[Mux.scala 31:69:@42206.4]
  assign _T_94394 = _T_94186 ? 16'h2 : _T_94393; // @[Mux.scala 31:69:@42207.4]
  assign _T_94395 = _T_94183 ? 16'h1 : _T_94394; // @[Mux.scala 31:69:@42208.4]
  assign _T_94396 = _T_94395[0]; // @[OneHot.scala 66:30:@42209.4]
  assign _T_94397 = _T_94395[1]; // @[OneHot.scala 66:30:@42210.4]
  assign _T_94398 = _T_94395[2]; // @[OneHot.scala 66:30:@42211.4]
  assign _T_94399 = _T_94395[3]; // @[OneHot.scala 66:30:@42212.4]
  assign _T_94400 = _T_94395[4]; // @[OneHot.scala 66:30:@42213.4]
  assign _T_94401 = _T_94395[5]; // @[OneHot.scala 66:30:@42214.4]
  assign _T_94402 = _T_94395[6]; // @[OneHot.scala 66:30:@42215.4]
  assign _T_94403 = _T_94395[7]; // @[OneHot.scala 66:30:@42216.4]
  assign _T_94404 = _T_94395[8]; // @[OneHot.scala 66:30:@42217.4]
  assign _T_94405 = _T_94395[9]; // @[OneHot.scala 66:30:@42218.4]
  assign _T_94406 = _T_94395[10]; // @[OneHot.scala 66:30:@42219.4]
  assign _T_94407 = _T_94395[11]; // @[OneHot.scala 66:30:@42220.4]
  assign _T_94408 = _T_94395[12]; // @[OneHot.scala 66:30:@42221.4]
  assign _T_94409 = _T_94395[13]; // @[OneHot.scala 66:30:@42222.4]
  assign _T_94410 = _T_94395[14]; // @[OneHot.scala 66:30:@42223.4]
  assign _T_94411 = _T_94395[15]; // @[OneHot.scala 66:30:@42224.4]
  assign _T_94452 = _T_94183 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42242.4]
  assign _T_94453 = _T_94180 ? 16'h4000 : _T_94452; // @[Mux.scala 31:69:@42243.4]
  assign _T_94454 = _T_94225 ? 16'h2000 : _T_94453; // @[Mux.scala 31:69:@42244.4]
  assign _T_94455 = _T_94222 ? 16'h1000 : _T_94454; // @[Mux.scala 31:69:@42245.4]
  assign _T_94456 = _T_94219 ? 16'h800 : _T_94455; // @[Mux.scala 31:69:@42246.4]
  assign _T_94457 = _T_94216 ? 16'h400 : _T_94456; // @[Mux.scala 31:69:@42247.4]
  assign _T_94458 = _T_94213 ? 16'h200 : _T_94457; // @[Mux.scala 31:69:@42248.4]
  assign _T_94459 = _T_94210 ? 16'h100 : _T_94458; // @[Mux.scala 31:69:@42249.4]
  assign _T_94460 = _T_94207 ? 16'h80 : _T_94459; // @[Mux.scala 31:69:@42250.4]
  assign _T_94461 = _T_94204 ? 16'h40 : _T_94460; // @[Mux.scala 31:69:@42251.4]
  assign _T_94462 = _T_94201 ? 16'h20 : _T_94461; // @[Mux.scala 31:69:@42252.4]
  assign _T_94463 = _T_94198 ? 16'h10 : _T_94462; // @[Mux.scala 31:69:@42253.4]
  assign _T_94464 = _T_94195 ? 16'h8 : _T_94463; // @[Mux.scala 31:69:@42254.4]
  assign _T_94465 = _T_94192 ? 16'h4 : _T_94464; // @[Mux.scala 31:69:@42255.4]
  assign _T_94466 = _T_94189 ? 16'h2 : _T_94465; // @[Mux.scala 31:69:@42256.4]
  assign _T_94467 = _T_94186 ? 16'h1 : _T_94466; // @[Mux.scala 31:69:@42257.4]
  assign _T_94468 = _T_94467[0]; // @[OneHot.scala 66:30:@42258.4]
  assign _T_94469 = _T_94467[1]; // @[OneHot.scala 66:30:@42259.4]
  assign _T_94470 = _T_94467[2]; // @[OneHot.scala 66:30:@42260.4]
  assign _T_94471 = _T_94467[3]; // @[OneHot.scala 66:30:@42261.4]
  assign _T_94472 = _T_94467[4]; // @[OneHot.scala 66:30:@42262.4]
  assign _T_94473 = _T_94467[5]; // @[OneHot.scala 66:30:@42263.4]
  assign _T_94474 = _T_94467[6]; // @[OneHot.scala 66:30:@42264.4]
  assign _T_94475 = _T_94467[7]; // @[OneHot.scala 66:30:@42265.4]
  assign _T_94476 = _T_94467[8]; // @[OneHot.scala 66:30:@42266.4]
  assign _T_94477 = _T_94467[9]; // @[OneHot.scala 66:30:@42267.4]
  assign _T_94478 = _T_94467[10]; // @[OneHot.scala 66:30:@42268.4]
  assign _T_94479 = _T_94467[11]; // @[OneHot.scala 66:30:@42269.4]
  assign _T_94480 = _T_94467[12]; // @[OneHot.scala 66:30:@42270.4]
  assign _T_94481 = _T_94467[13]; // @[OneHot.scala 66:30:@42271.4]
  assign _T_94482 = _T_94467[14]; // @[OneHot.scala 66:30:@42272.4]
  assign _T_94483 = _T_94467[15]; // @[OneHot.scala 66:30:@42273.4]
  assign _T_94524 = _T_94186 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42291.4]
  assign _T_94525 = _T_94183 ? 16'h4000 : _T_94524; // @[Mux.scala 31:69:@42292.4]
  assign _T_94526 = _T_94180 ? 16'h2000 : _T_94525; // @[Mux.scala 31:69:@42293.4]
  assign _T_94527 = _T_94225 ? 16'h1000 : _T_94526; // @[Mux.scala 31:69:@42294.4]
  assign _T_94528 = _T_94222 ? 16'h800 : _T_94527; // @[Mux.scala 31:69:@42295.4]
  assign _T_94529 = _T_94219 ? 16'h400 : _T_94528; // @[Mux.scala 31:69:@42296.4]
  assign _T_94530 = _T_94216 ? 16'h200 : _T_94529; // @[Mux.scala 31:69:@42297.4]
  assign _T_94531 = _T_94213 ? 16'h100 : _T_94530; // @[Mux.scala 31:69:@42298.4]
  assign _T_94532 = _T_94210 ? 16'h80 : _T_94531; // @[Mux.scala 31:69:@42299.4]
  assign _T_94533 = _T_94207 ? 16'h40 : _T_94532; // @[Mux.scala 31:69:@42300.4]
  assign _T_94534 = _T_94204 ? 16'h20 : _T_94533; // @[Mux.scala 31:69:@42301.4]
  assign _T_94535 = _T_94201 ? 16'h10 : _T_94534; // @[Mux.scala 31:69:@42302.4]
  assign _T_94536 = _T_94198 ? 16'h8 : _T_94535; // @[Mux.scala 31:69:@42303.4]
  assign _T_94537 = _T_94195 ? 16'h4 : _T_94536; // @[Mux.scala 31:69:@42304.4]
  assign _T_94538 = _T_94192 ? 16'h2 : _T_94537; // @[Mux.scala 31:69:@42305.4]
  assign _T_94539 = _T_94189 ? 16'h1 : _T_94538; // @[Mux.scala 31:69:@42306.4]
  assign _T_94540 = _T_94539[0]; // @[OneHot.scala 66:30:@42307.4]
  assign _T_94541 = _T_94539[1]; // @[OneHot.scala 66:30:@42308.4]
  assign _T_94542 = _T_94539[2]; // @[OneHot.scala 66:30:@42309.4]
  assign _T_94543 = _T_94539[3]; // @[OneHot.scala 66:30:@42310.4]
  assign _T_94544 = _T_94539[4]; // @[OneHot.scala 66:30:@42311.4]
  assign _T_94545 = _T_94539[5]; // @[OneHot.scala 66:30:@42312.4]
  assign _T_94546 = _T_94539[6]; // @[OneHot.scala 66:30:@42313.4]
  assign _T_94547 = _T_94539[7]; // @[OneHot.scala 66:30:@42314.4]
  assign _T_94548 = _T_94539[8]; // @[OneHot.scala 66:30:@42315.4]
  assign _T_94549 = _T_94539[9]; // @[OneHot.scala 66:30:@42316.4]
  assign _T_94550 = _T_94539[10]; // @[OneHot.scala 66:30:@42317.4]
  assign _T_94551 = _T_94539[11]; // @[OneHot.scala 66:30:@42318.4]
  assign _T_94552 = _T_94539[12]; // @[OneHot.scala 66:30:@42319.4]
  assign _T_94553 = _T_94539[13]; // @[OneHot.scala 66:30:@42320.4]
  assign _T_94554 = _T_94539[14]; // @[OneHot.scala 66:30:@42321.4]
  assign _T_94555 = _T_94539[15]; // @[OneHot.scala 66:30:@42322.4]
  assign _T_94596 = _T_94189 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42340.4]
  assign _T_94597 = _T_94186 ? 16'h4000 : _T_94596; // @[Mux.scala 31:69:@42341.4]
  assign _T_94598 = _T_94183 ? 16'h2000 : _T_94597; // @[Mux.scala 31:69:@42342.4]
  assign _T_94599 = _T_94180 ? 16'h1000 : _T_94598; // @[Mux.scala 31:69:@42343.4]
  assign _T_94600 = _T_94225 ? 16'h800 : _T_94599; // @[Mux.scala 31:69:@42344.4]
  assign _T_94601 = _T_94222 ? 16'h400 : _T_94600; // @[Mux.scala 31:69:@42345.4]
  assign _T_94602 = _T_94219 ? 16'h200 : _T_94601; // @[Mux.scala 31:69:@42346.4]
  assign _T_94603 = _T_94216 ? 16'h100 : _T_94602; // @[Mux.scala 31:69:@42347.4]
  assign _T_94604 = _T_94213 ? 16'h80 : _T_94603; // @[Mux.scala 31:69:@42348.4]
  assign _T_94605 = _T_94210 ? 16'h40 : _T_94604; // @[Mux.scala 31:69:@42349.4]
  assign _T_94606 = _T_94207 ? 16'h20 : _T_94605; // @[Mux.scala 31:69:@42350.4]
  assign _T_94607 = _T_94204 ? 16'h10 : _T_94606; // @[Mux.scala 31:69:@42351.4]
  assign _T_94608 = _T_94201 ? 16'h8 : _T_94607; // @[Mux.scala 31:69:@42352.4]
  assign _T_94609 = _T_94198 ? 16'h4 : _T_94608; // @[Mux.scala 31:69:@42353.4]
  assign _T_94610 = _T_94195 ? 16'h2 : _T_94609; // @[Mux.scala 31:69:@42354.4]
  assign _T_94611 = _T_94192 ? 16'h1 : _T_94610; // @[Mux.scala 31:69:@42355.4]
  assign _T_94612 = _T_94611[0]; // @[OneHot.scala 66:30:@42356.4]
  assign _T_94613 = _T_94611[1]; // @[OneHot.scala 66:30:@42357.4]
  assign _T_94614 = _T_94611[2]; // @[OneHot.scala 66:30:@42358.4]
  assign _T_94615 = _T_94611[3]; // @[OneHot.scala 66:30:@42359.4]
  assign _T_94616 = _T_94611[4]; // @[OneHot.scala 66:30:@42360.4]
  assign _T_94617 = _T_94611[5]; // @[OneHot.scala 66:30:@42361.4]
  assign _T_94618 = _T_94611[6]; // @[OneHot.scala 66:30:@42362.4]
  assign _T_94619 = _T_94611[7]; // @[OneHot.scala 66:30:@42363.4]
  assign _T_94620 = _T_94611[8]; // @[OneHot.scala 66:30:@42364.4]
  assign _T_94621 = _T_94611[9]; // @[OneHot.scala 66:30:@42365.4]
  assign _T_94622 = _T_94611[10]; // @[OneHot.scala 66:30:@42366.4]
  assign _T_94623 = _T_94611[11]; // @[OneHot.scala 66:30:@42367.4]
  assign _T_94624 = _T_94611[12]; // @[OneHot.scala 66:30:@42368.4]
  assign _T_94625 = _T_94611[13]; // @[OneHot.scala 66:30:@42369.4]
  assign _T_94626 = _T_94611[14]; // @[OneHot.scala 66:30:@42370.4]
  assign _T_94627 = _T_94611[15]; // @[OneHot.scala 66:30:@42371.4]
  assign _T_94668 = _T_94192 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42389.4]
  assign _T_94669 = _T_94189 ? 16'h4000 : _T_94668; // @[Mux.scala 31:69:@42390.4]
  assign _T_94670 = _T_94186 ? 16'h2000 : _T_94669; // @[Mux.scala 31:69:@42391.4]
  assign _T_94671 = _T_94183 ? 16'h1000 : _T_94670; // @[Mux.scala 31:69:@42392.4]
  assign _T_94672 = _T_94180 ? 16'h800 : _T_94671; // @[Mux.scala 31:69:@42393.4]
  assign _T_94673 = _T_94225 ? 16'h400 : _T_94672; // @[Mux.scala 31:69:@42394.4]
  assign _T_94674 = _T_94222 ? 16'h200 : _T_94673; // @[Mux.scala 31:69:@42395.4]
  assign _T_94675 = _T_94219 ? 16'h100 : _T_94674; // @[Mux.scala 31:69:@42396.4]
  assign _T_94676 = _T_94216 ? 16'h80 : _T_94675; // @[Mux.scala 31:69:@42397.4]
  assign _T_94677 = _T_94213 ? 16'h40 : _T_94676; // @[Mux.scala 31:69:@42398.4]
  assign _T_94678 = _T_94210 ? 16'h20 : _T_94677; // @[Mux.scala 31:69:@42399.4]
  assign _T_94679 = _T_94207 ? 16'h10 : _T_94678; // @[Mux.scala 31:69:@42400.4]
  assign _T_94680 = _T_94204 ? 16'h8 : _T_94679; // @[Mux.scala 31:69:@42401.4]
  assign _T_94681 = _T_94201 ? 16'h4 : _T_94680; // @[Mux.scala 31:69:@42402.4]
  assign _T_94682 = _T_94198 ? 16'h2 : _T_94681; // @[Mux.scala 31:69:@42403.4]
  assign _T_94683 = _T_94195 ? 16'h1 : _T_94682; // @[Mux.scala 31:69:@42404.4]
  assign _T_94684 = _T_94683[0]; // @[OneHot.scala 66:30:@42405.4]
  assign _T_94685 = _T_94683[1]; // @[OneHot.scala 66:30:@42406.4]
  assign _T_94686 = _T_94683[2]; // @[OneHot.scala 66:30:@42407.4]
  assign _T_94687 = _T_94683[3]; // @[OneHot.scala 66:30:@42408.4]
  assign _T_94688 = _T_94683[4]; // @[OneHot.scala 66:30:@42409.4]
  assign _T_94689 = _T_94683[5]; // @[OneHot.scala 66:30:@42410.4]
  assign _T_94690 = _T_94683[6]; // @[OneHot.scala 66:30:@42411.4]
  assign _T_94691 = _T_94683[7]; // @[OneHot.scala 66:30:@42412.4]
  assign _T_94692 = _T_94683[8]; // @[OneHot.scala 66:30:@42413.4]
  assign _T_94693 = _T_94683[9]; // @[OneHot.scala 66:30:@42414.4]
  assign _T_94694 = _T_94683[10]; // @[OneHot.scala 66:30:@42415.4]
  assign _T_94695 = _T_94683[11]; // @[OneHot.scala 66:30:@42416.4]
  assign _T_94696 = _T_94683[12]; // @[OneHot.scala 66:30:@42417.4]
  assign _T_94697 = _T_94683[13]; // @[OneHot.scala 66:30:@42418.4]
  assign _T_94698 = _T_94683[14]; // @[OneHot.scala 66:30:@42419.4]
  assign _T_94699 = _T_94683[15]; // @[OneHot.scala 66:30:@42420.4]
  assign _T_94740 = _T_94195 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42438.4]
  assign _T_94741 = _T_94192 ? 16'h4000 : _T_94740; // @[Mux.scala 31:69:@42439.4]
  assign _T_94742 = _T_94189 ? 16'h2000 : _T_94741; // @[Mux.scala 31:69:@42440.4]
  assign _T_94743 = _T_94186 ? 16'h1000 : _T_94742; // @[Mux.scala 31:69:@42441.4]
  assign _T_94744 = _T_94183 ? 16'h800 : _T_94743; // @[Mux.scala 31:69:@42442.4]
  assign _T_94745 = _T_94180 ? 16'h400 : _T_94744; // @[Mux.scala 31:69:@42443.4]
  assign _T_94746 = _T_94225 ? 16'h200 : _T_94745; // @[Mux.scala 31:69:@42444.4]
  assign _T_94747 = _T_94222 ? 16'h100 : _T_94746; // @[Mux.scala 31:69:@42445.4]
  assign _T_94748 = _T_94219 ? 16'h80 : _T_94747; // @[Mux.scala 31:69:@42446.4]
  assign _T_94749 = _T_94216 ? 16'h40 : _T_94748; // @[Mux.scala 31:69:@42447.4]
  assign _T_94750 = _T_94213 ? 16'h20 : _T_94749; // @[Mux.scala 31:69:@42448.4]
  assign _T_94751 = _T_94210 ? 16'h10 : _T_94750; // @[Mux.scala 31:69:@42449.4]
  assign _T_94752 = _T_94207 ? 16'h8 : _T_94751; // @[Mux.scala 31:69:@42450.4]
  assign _T_94753 = _T_94204 ? 16'h4 : _T_94752; // @[Mux.scala 31:69:@42451.4]
  assign _T_94754 = _T_94201 ? 16'h2 : _T_94753; // @[Mux.scala 31:69:@42452.4]
  assign _T_94755 = _T_94198 ? 16'h1 : _T_94754; // @[Mux.scala 31:69:@42453.4]
  assign _T_94756 = _T_94755[0]; // @[OneHot.scala 66:30:@42454.4]
  assign _T_94757 = _T_94755[1]; // @[OneHot.scala 66:30:@42455.4]
  assign _T_94758 = _T_94755[2]; // @[OneHot.scala 66:30:@42456.4]
  assign _T_94759 = _T_94755[3]; // @[OneHot.scala 66:30:@42457.4]
  assign _T_94760 = _T_94755[4]; // @[OneHot.scala 66:30:@42458.4]
  assign _T_94761 = _T_94755[5]; // @[OneHot.scala 66:30:@42459.4]
  assign _T_94762 = _T_94755[6]; // @[OneHot.scala 66:30:@42460.4]
  assign _T_94763 = _T_94755[7]; // @[OneHot.scala 66:30:@42461.4]
  assign _T_94764 = _T_94755[8]; // @[OneHot.scala 66:30:@42462.4]
  assign _T_94765 = _T_94755[9]; // @[OneHot.scala 66:30:@42463.4]
  assign _T_94766 = _T_94755[10]; // @[OneHot.scala 66:30:@42464.4]
  assign _T_94767 = _T_94755[11]; // @[OneHot.scala 66:30:@42465.4]
  assign _T_94768 = _T_94755[12]; // @[OneHot.scala 66:30:@42466.4]
  assign _T_94769 = _T_94755[13]; // @[OneHot.scala 66:30:@42467.4]
  assign _T_94770 = _T_94755[14]; // @[OneHot.scala 66:30:@42468.4]
  assign _T_94771 = _T_94755[15]; // @[OneHot.scala 66:30:@42469.4]
  assign _T_94812 = _T_94198 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42487.4]
  assign _T_94813 = _T_94195 ? 16'h4000 : _T_94812; // @[Mux.scala 31:69:@42488.4]
  assign _T_94814 = _T_94192 ? 16'h2000 : _T_94813; // @[Mux.scala 31:69:@42489.4]
  assign _T_94815 = _T_94189 ? 16'h1000 : _T_94814; // @[Mux.scala 31:69:@42490.4]
  assign _T_94816 = _T_94186 ? 16'h800 : _T_94815; // @[Mux.scala 31:69:@42491.4]
  assign _T_94817 = _T_94183 ? 16'h400 : _T_94816; // @[Mux.scala 31:69:@42492.4]
  assign _T_94818 = _T_94180 ? 16'h200 : _T_94817; // @[Mux.scala 31:69:@42493.4]
  assign _T_94819 = _T_94225 ? 16'h100 : _T_94818; // @[Mux.scala 31:69:@42494.4]
  assign _T_94820 = _T_94222 ? 16'h80 : _T_94819; // @[Mux.scala 31:69:@42495.4]
  assign _T_94821 = _T_94219 ? 16'h40 : _T_94820; // @[Mux.scala 31:69:@42496.4]
  assign _T_94822 = _T_94216 ? 16'h20 : _T_94821; // @[Mux.scala 31:69:@42497.4]
  assign _T_94823 = _T_94213 ? 16'h10 : _T_94822; // @[Mux.scala 31:69:@42498.4]
  assign _T_94824 = _T_94210 ? 16'h8 : _T_94823; // @[Mux.scala 31:69:@42499.4]
  assign _T_94825 = _T_94207 ? 16'h4 : _T_94824; // @[Mux.scala 31:69:@42500.4]
  assign _T_94826 = _T_94204 ? 16'h2 : _T_94825; // @[Mux.scala 31:69:@42501.4]
  assign _T_94827 = _T_94201 ? 16'h1 : _T_94826; // @[Mux.scala 31:69:@42502.4]
  assign _T_94828 = _T_94827[0]; // @[OneHot.scala 66:30:@42503.4]
  assign _T_94829 = _T_94827[1]; // @[OneHot.scala 66:30:@42504.4]
  assign _T_94830 = _T_94827[2]; // @[OneHot.scala 66:30:@42505.4]
  assign _T_94831 = _T_94827[3]; // @[OneHot.scala 66:30:@42506.4]
  assign _T_94832 = _T_94827[4]; // @[OneHot.scala 66:30:@42507.4]
  assign _T_94833 = _T_94827[5]; // @[OneHot.scala 66:30:@42508.4]
  assign _T_94834 = _T_94827[6]; // @[OneHot.scala 66:30:@42509.4]
  assign _T_94835 = _T_94827[7]; // @[OneHot.scala 66:30:@42510.4]
  assign _T_94836 = _T_94827[8]; // @[OneHot.scala 66:30:@42511.4]
  assign _T_94837 = _T_94827[9]; // @[OneHot.scala 66:30:@42512.4]
  assign _T_94838 = _T_94827[10]; // @[OneHot.scala 66:30:@42513.4]
  assign _T_94839 = _T_94827[11]; // @[OneHot.scala 66:30:@42514.4]
  assign _T_94840 = _T_94827[12]; // @[OneHot.scala 66:30:@42515.4]
  assign _T_94841 = _T_94827[13]; // @[OneHot.scala 66:30:@42516.4]
  assign _T_94842 = _T_94827[14]; // @[OneHot.scala 66:30:@42517.4]
  assign _T_94843 = _T_94827[15]; // @[OneHot.scala 66:30:@42518.4]
  assign _T_94884 = _T_94201 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42536.4]
  assign _T_94885 = _T_94198 ? 16'h4000 : _T_94884; // @[Mux.scala 31:69:@42537.4]
  assign _T_94886 = _T_94195 ? 16'h2000 : _T_94885; // @[Mux.scala 31:69:@42538.4]
  assign _T_94887 = _T_94192 ? 16'h1000 : _T_94886; // @[Mux.scala 31:69:@42539.4]
  assign _T_94888 = _T_94189 ? 16'h800 : _T_94887; // @[Mux.scala 31:69:@42540.4]
  assign _T_94889 = _T_94186 ? 16'h400 : _T_94888; // @[Mux.scala 31:69:@42541.4]
  assign _T_94890 = _T_94183 ? 16'h200 : _T_94889; // @[Mux.scala 31:69:@42542.4]
  assign _T_94891 = _T_94180 ? 16'h100 : _T_94890; // @[Mux.scala 31:69:@42543.4]
  assign _T_94892 = _T_94225 ? 16'h80 : _T_94891; // @[Mux.scala 31:69:@42544.4]
  assign _T_94893 = _T_94222 ? 16'h40 : _T_94892; // @[Mux.scala 31:69:@42545.4]
  assign _T_94894 = _T_94219 ? 16'h20 : _T_94893; // @[Mux.scala 31:69:@42546.4]
  assign _T_94895 = _T_94216 ? 16'h10 : _T_94894; // @[Mux.scala 31:69:@42547.4]
  assign _T_94896 = _T_94213 ? 16'h8 : _T_94895; // @[Mux.scala 31:69:@42548.4]
  assign _T_94897 = _T_94210 ? 16'h4 : _T_94896; // @[Mux.scala 31:69:@42549.4]
  assign _T_94898 = _T_94207 ? 16'h2 : _T_94897; // @[Mux.scala 31:69:@42550.4]
  assign _T_94899 = _T_94204 ? 16'h1 : _T_94898; // @[Mux.scala 31:69:@42551.4]
  assign _T_94900 = _T_94899[0]; // @[OneHot.scala 66:30:@42552.4]
  assign _T_94901 = _T_94899[1]; // @[OneHot.scala 66:30:@42553.4]
  assign _T_94902 = _T_94899[2]; // @[OneHot.scala 66:30:@42554.4]
  assign _T_94903 = _T_94899[3]; // @[OneHot.scala 66:30:@42555.4]
  assign _T_94904 = _T_94899[4]; // @[OneHot.scala 66:30:@42556.4]
  assign _T_94905 = _T_94899[5]; // @[OneHot.scala 66:30:@42557.4]
  assign _T_94906 = _T_94899[6]; // @[OneHot.scala 66:30:@42558.4]
  assign _T_94907 = _T_94899[7]; // @[OneHot.scala 66:30:@42559.4]
  assign _T_94908 = _T_94899[8]; // @[OneHot.scala 66:30:@42560.4]
  assign _T_94909 = _T_94899[9]; // @[OneHot.scala 66:30:@42561.4]
  assign _T_94910 = _T_94899[10]; // @[OneHot.scala 66:30:@42562.4]
  assign _T_94911 = _T_94899[11]; // @[OneHot.scala 66:30:@42563.4]
  assign _T_94912 = _T_94899[12]; // @[OneHot.scala 66:30:@42564.4]
  assign _T_94913 = _T_94899[13]; // @[OneHot.scala 66:30:@42565.4]
  assign _T_94914 = _T_94899[14]; // @[OneHot.scala 66:30:@42566.4]
  assign _T_94915 = _T_94899[15]; // @[OneHot.scala 66:30:@42567.4]
  assign _T_94956 = _T_94204 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42585.4]
  assign _T_94957 = _T_94201 ? 16'h4000 : _T_94956; // @[Mux.scala 31:69:@42586.4]
  assign _T_94958 = _T_94198 ? 16'h2000 : _T_94957; // @[Mux.scala 31:69:@42587.4]
  assign _T_94959 = _T_94195 ? 16'h1000 : _T_94958; // @[Mux.scala 31:69:@42588.4]
  assign _T_94960 = _T_94192 ? 16'h800 : _T_94959; // @[Mux.scala 31:69:@42589.4]
  assign _T_94961 = _T_94189 ? 16'h400 : _T_94960; // @[Mux.scala 31:69:@42590.4]
  assign _T_94962 = _T_94186 ? 16'h200 : _T_94961; // @[Mux.scala 31:69:@42591.4]
  assign _T_94963 = _T_94183 ? 16'h100 : _T_94962; // @[Mux.scala 31:69:@42592.4]
  assign _T_94964 = _T_94180 ? 16'h80 : _T_94963; // @[Mux.scala 31:69:@42593.4]
  assign _T_94965 = _T_94225 ? 16'h40 : _T_94964; // @[Mux.scala 31:69:@42594.4]
  assign _T_94966 = _T_94222 ? 16'h20 : _T_94965; // @[Mux.scala 31:69:@42595.4]
  assign _T_94967 = _T_94219 ? 16'h10 : _T_94966; // @[Mux.scala 31:69:@42596.4]
  assign _T_94968 = _T_94216 ? 16'h8 : _T_94967; // @[Mux.scala 31:69:@42597.4]
  assign _T_94969 = _T_94213 ? 16'h4 : _T_94968; // @[Mux.scala 31:69:@42598.4]
  assign _T_94970 = _T_94210 ? 16'h2 : _T_94969; // @[Mux.scala 31:69:@42599.4]
  assign _T_94971 = _T_94207 ? 16'h1 : _T_94970; // @[Mux.scala 31:69:@42600.4]
  assign _T_94972 = _T_94971[0]; // @[OneHot.scala 66:30:@42601.4]
  assign _T_94973 = _T_94971[1]; // @[OneHot.scala 66:30:@42602.4]
  assign _T_94974 = _T_94971[2]; // @[OneHot.scala 66:30:@42603.4]
  assign _T_94975 = _T_94971[3]; // @[OneHot.scala 66:30:@42604.4]
  assign _T_94976 = _T_94971[4]; // @[OneHot.scala 66:30:@42605.4]
  assign _T_94977 = _T_94971[5]; // @[OneHot.scala 66:30:@42606.4]
  assign _T_94978 = _T_94971[6]; // @[OneHot.scala 66:30:@42607.4]
  assign _T_94979 = _T_94971[7]; // @[OneHot.scala 66:30:@42608.4]
  assign _T_94980 = _T_94971[8]; // @[OneHot.scala 66:30:@42609.4]
  assign _T_94981 = _T_94971[9]; // @[OneHot.scala 66:30:@42610.4]
  assign _T_94982 = _T_94971[10]; // @[OneHot.scala 66:30:@42611.4]
  assign _T_94983 = _T_94971[11]; // @[OneHot.scala 66:30:@42612.4]
  assign _T_94984 = _T_94971[12]; // @[OneHot.scala 66:30:@42613.4]
  assign _T_94985 = _T_94971[13]; // @[OneHot.scala 66:30:@42614.4]
  assign _T_94986 = _T_94971[14]; // @[OneHot.scala 66:30:@42615.4]
  assign _T_94987 = _T_94971[15]; // @[OneHot.scala 66:30:@42616.4]
  assign _T_95028 = _T_94207 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42634.4]
  assign _T_95029 = _T_94204 ? 16'h4000 : _T_95028; // @[Mux.scala 31:69:@42635.4]
  assign _T_95030 = _T_94201 ? 16'h2000 : _T_95029; // @[Mux.scala 31:69:@42636.4]
  assign _T_95031 = _T_94198 ? 16'h1000 : _T_95030; // @[Mux.scala 31:69:@42637.4]
  assign _T_95032 = _T_94195 ? 16'h800 : _T_95031; // @[Mux.scala 31:69:@42638.4]
  assign _T_95033 = _T_94192 ? 16'h400 : _T_95032; // @[Mux.scala 31:69:@42639.4]
  assign _T_95034 = _T_94189 ? 16'h200 : _T_95033; // @[Mux.scala 31:69:@42640.4]
  assign _T_95035 = _T_94186 ? 16'h100 : _T_95034; // @[Mux.scala 31:69:@42641.4]
  assign _T_95036 = _T_94183 ? 16'h80 : _T_95035; // @[Mux.scala 31:69:@42642.4]
  assign _T_95037 = _T_94180 ? 16'h40 : _T_95036; // @[Mux.scala 31:69:@42643.4]
  assign _T_95038 = _T_94225 ? 16'h20 : _T_95037; // @[Mux.scala 31:69:@42644.4]
  assign _T_95039 = _T_94222 ? 16'h10 : _T_95038; // @[Mux.scala 31:69:@42645.4]
  assign _T_95040 = _T_94219 ? 16'h8 : _T_95039; // @[Mux.scala 31:69:@42646.4]
  assign _T_95041 = _T_94216 ? 16'h4 : _T_95040; // @[Mux.scala 31:69:@42647.4]
  assign _T_95042 = _T_94213 ? 16'h2 : _T_95041; // @[Mux.scala 31:69:@42648.4]
  assign _T_95043 = _T_94210 ? 16'h1 : _T_95042; // @[Mux.scala 31:69:@42649.4]
  assign _T_95044 = _T_95043[0]; // @[OneHot.scala 66:30:@42650.4]
  assign _T_95045 = _T_95043[1]; // @[OneHot.scala 66:30:@42651.4]
  assign _T_95046 = _T_95043[2]; // @[OneHot.scala 66:30:@42652.4]
  assign _T_95047 = _T_95043[3]; // @[OneHot.scala 66:30:@42653.4]
  assign _T_95048 = _T_95043[4]; // @[OneHot.scala 66:30:@42654.4]
  assign _T_95049 = _T_95043[5]; // @[OneHot.scala 66:30:@42655.4]
  assign _T_95050 = _T_95043[6]; // @[OneHot.scala 66:30:@42656.4]
  assign _T_95051 = _T_95043[7]; // @[OneHot.scala 66:30:@42657.4]
  assign _T_95052 = _T_95043[8]; // @[OneHot.scala 66:30:@42658.4]
  assign _T_95053 = _T_95043[9]; // @[OneHot.scala 66:30:@42659.4]
  assign _T_95054 = _T_95043[10]; // @[OneHot.scala 66:30:@42660.4]
  assign _T_95055 = _T_95043[11]; // @[OneHot.scala 66:30:@42661.4]
  assign _T_95056 = _T_95043[12]; // @[OneHot.scala 66:30:@42662.4]
  assign _T_95057 = _T_95043[13]; // @[OneHot.scala 66:30:@42663.4]
  assign _T_95058 = _T_95043[14]; // @[OneHot.scala 66:30:@42664.4]
  assign _T_95059 = _T_95043[15]; // @[OneHot.scala 66:30:@42665.4]
  assign _T_95100 = _T_94210 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42683.4]
  assign _T_95101 = _T_94207 ? 16'h4000 : _T_95100; // @[Mux.scala 31:69:@42684.4]
  assign _T_95102 = _T_94204 ? 16'h2000 : _T_95101; // @[Mux.scala 31:69:@42685.4]
  assign _T_95103 = _T_94201 ? 16'h1000 : _T_95102; // @[Mux.scala 31:69:@42686.4]
  assign _T_95104 = _T_94198 ? 16'h800 : _T_95103; // @[Mux.scala 31:69:@42687.4]
  assign _T_95105 = _T_94195 ? 16'h400 : _T_95104; // @[Mux.scala 31:69:@42688.4]
  assign _T_95106 = _T_94192 ? 16'h200 : _T_95105; // @[Mux.scala 31:69:@42689.4]
  assign _T_95107 = _T_94189 ? 16'h100 : _T_95106; // @[Mux.scala 31:69:@42690.4]
  assign _T_95108 = _T_94186 ? 16'h80 : _T_95107; // @[Mux.scala 31:69:@42691.4]
  assign _T_95109 = _T_94183 ? 16'h40 : _T_95108; // @[Mux.scala 31:69:@42692.4]
  assign _T_95110 = _T_94180 ? 16'h20 : _T_95109; // @[Mux.scala 31:69:@42693.4]
  assign _T_95111 = _T_94225 ? 16'h10 : _T_95110; // @[Mux.scala 31:69:@42694.4]
  assign _T_95112 = _T_94222 ? 16'h8 : _T_95111; // @[Mux.scala 31:69:@42695.4]
  assign _T_95113 = _T_94219 ? 16'h4 : _T_95112; // @[Mux.scala 31:69:@42696.4]
  assign _T_95114 = _T_94216 ? 16'h2 : _T_95113; // @[Mux.scala 31:69:@42697.4]
  assign _T_95115 = _T_94213 ? 16'h1 : _T_95114; // @[Mux.scala 31:69:@42698.4]
  assign _T_95116 = _T_95115[0]; // @[OneHot.scala 66:30:@42699.4]
  assign _T_95117 = _T_95115[1]; // @[OneHot.scala 66:30:@42700.4]
  assign _T_95118 = _T_95115[2]; // @[OneHot.scala 66:30:@42701.4]
  assign _T_95119 = _T_95115[3]; // @[OneHot.scala 66:30:@42702.4]
  assign _T_95120 = _T_95115[4]; // @[OneHot.scala 66:30:@42703.4]
  assign _T_95121 = _T_95115[5]; // @[OneHot.scala 66:30:@42704.4]
  assign _T_95122 = _T_95115[6]; // @[OneHot.scala 66:30:@42705.4]
  assign _T_95123 = _T_95115[7]; // @[OneHot.scala 66:30:@42706.4]
  assign _T_95124 = _T_95115[8]; // @[OneHot.scala 66:30:@42707.4]
  assign _T_95125 = _T_95115[9]; // @[OneHot.scala 66:30:@42708.4]
  assign _T_95126 = _T_95115[10]; // @[OneHot.scala 66:30:@42709.4]
  assign _T_95127 = _T_95115[11]; // @[OneHot.scala 66:30:@42710.4]
  assign _T_95128 = _T_95115[12]; // @[OneHot.scala 66:30:@42711.4]
  assign _T_95129 = _T_95115[13]; // @[OneHot.scala 66:30:@42712.4]
  assign _T_95130 = _T_95115[14]; // @[OneHot.scala 66:30:@42713.4]
  assign _T_95131 = _T_95115[15]; // @[OneHot.scala 66:30:@42714.4]
  assign _T_95172 = _T_94213 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42732.4]
  assign _T_95173 = _T_94210 ? 16'h4000 : _T_95172; // @[Mux.scala 31:69:@42733.4]
  assign _T_95174 = _T_94207 ? 16'h2000 : _T_95173; // @[Mux.scala 31:69:@42734.4]
  assign _T_95175 = _T_94204 ? 16'h1000 : _T_95174; // @[Mux.scala 31:69:@42735.4]
  assign _T_95176 = _T_94201 ? 16'h800 : _T_95175; // @[Mux.scala 31:69:@42736.4]
  assign _T_95177 = _T_94198 ? 16'h400 : _T_95176; // @[Mux.scala 31:69:@42737.4]
  assign _T_95178 = _T_94195 ? 16'h200 : _T_95177; // @[Mux.scala 31:69:@42738.4]
  assign _T_95179 = _T_94192 ? 16'h100 : _T_95178; // @[Mux.scala 31:69:@42739.4]
  assign _T_95180 = _T_94189 ? 16'h80 : _T_95179; // @[Mux.scala 31:69:@42740.4]
  assign _T_95181 = _T_94186 ? 16'h40 : _T_95180; // @[Mux.scala 31:69:@42741.4]
  assign _T_95182 = _T_94183 ? 16'h20 : _T_95181; // @[Mux.scala 31:69:@42742.4]
  assign _T_95183 = _T_94180 ? 16'h10 : _T_95182; // @[Mux.scala 31:69:@42743.4]
  assign _T_95184 = _T_94225 ? 16'h8 : _T_95183; // @[Mux.scala 31:69:@42744.4]
  assign _T_95185 = _T_94222 ? 16'h4 : _T_95184; // @[Mux.scala 31:69:@42745.4]
  assign _T_95186 = _T_94219 ? 16'h2 : _T_95185; // @[Mux.scala 31:69:@42746.4]
  assign _T_95187 = _T_94216 ? 16'h1 : _T_95186; // @[Mux.scala 31:69:@42747.4]
  assign _T_95188 = _T_95187[0]; // @[OneHot.scala 66:30:@42748.4]
  assign _T_95189 = _T_95187[1]; // @[OneHot.scala 66:30:@42749.4]
  assign _T_95190 = _T_95187[2]; // @[OneHot.scala 66:30:@42750.4]
  assign _T_95191 = _T_95187[3]; // @[OneHot.scala 66:30:@42751.4]
  assign _T_95192 = _T_95187[4]; // @[OneHot.scala 66:30:@42752.4]
  assign _T_95193 = _T_95187[5]; // @[OneHot.scala 66:30:@42753.4]
  assign _T_95194 = _T_95187[6]; // @[OneHot.scala 66:30:@42754.4]
  assign _T_95195 = _T_95187[7]; // @[OneHot.scala 66:30:@42755.4]
  assign _T_95196 = _T_95187[8]; // @[OneHot.scala 66:30:@42756.4]
  assign _T_95197 = _T_95187[9]; // @[OneHot.scala 66:30:@42757.4]
  assign _T_95198 = _T_95187[10]; // @[OneHot.scala 66:30:@42758.4]
  assign _T_95199 = _T_95187[11]; // @[OneHot.scala 66:30:@42759.4]
  assign _T_95200 = _T_95187[12]; // @[OneHot.scala 66:30:@42760.4]
  assign _T_95201 = _T_95187[13]; // @[OneHot.scala 66:30:@42761.4]
  assign _T_95202 = _T_95187[14]; // @[OneHot.scala 66:30:@42762.4]
  assign _T_95203 = _T_95187[15]; // @[OneHot.scala 66:30:@42763.4]
  assign _T_95244 = _T_94216 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42781.4]
  assign _T_95245 = _T_94213 ? 16'h4000 : _T_95244; // @[Mux.scala 31:69:@42782.4]
  assign _T_95246 = _T_94210 ? 16'h2000 : _T_95245; // @[Mux.scala 31:69:@42783.4]
  assign _T_95247 = _T_94207 ? 16'h1000 : _T_95246; // @[Mux.scala 31:69:@42784.4]
  assign _T_95248 = _T_94204 ? 16'h800 : _T_95247; // @[Mux.scala 31:69:@42785.4]
  assign _T_95249 = _T_94201 ? 16'h400 : _T_95248; // @[Mux.scala 31:69:@42786.4]
  assign _T_95250 = _T_94198 ? 16'h200 : _T_95249; // @[Mux.scala 31:69:@42787.4]
  assign _T_95251 = _T_94195 ? 16'h100 : _T_95250; // @[Mux.scala 31:69:@42788.4]
  assign _T_95252 = _T_94192 ? 16'h80 : _T_95251; // @[Mux.scala 31:69:@42789.4]
  assign _T_95253 = _T_94189 ? 16'h40 : _T_95252; // @[Mux.scala 31:69:@42790.4]
  assign _T_95254 = _T_94186 ? 16'h20 : _T_95253; // @[Mux.scala 31:69:@42791.4]
  assign _T_95255 = _T_94183 ? 16'h10 : _T_95254; // @[Mux.scala 31:69:@42792.4]
  assign _T_95256 = _T_94180 ? 16'h8 : _T_95255; // @[Mux.scala 31:69:@42793.4]
  assign _T_95257 = _T_94225 ? 16'h4 : _T_95256; // @[Mux.scala 31:69:@42794.4]
  assign _T_95258 = _T_94222 ? 16'h2 : _T_95257; // @[Mux.scala 31:69:@42795.4]
  assign _T_95259 = _T_94219 ? 16'h1 : _T_95258; // @[Mux.scala 31:69:@42796.4]
  assign _T_95260 = _T_95259[0]; // @[OneHot.scala 66:30:@42797.4]
  assign _T_95261 = _T_95259[1]; // @[OneHot.scala 66:30:@42798.4]
  assign _T_95262 = _T_95259[2]; // @[OneHot.scala 66:30:@42799.4]
  assign _T_95263 = _T_95259[3]; // @[OneHot.scala 66:30:@42800.4]
  assign _T_95264 = _T_95259[4]; // @[OneHot.scala 66:30:@42801.4]
  assign _T_95265 = _T_95259[5]; // @[OneHot.scala 66:30:@42802.4]
  assign _T_95266 = _T_95259[6]; // @[OneHot.scala 66:30:@42803.4]
  assign _T_95267 = _T_95259[7]; // @[OneHot.scala 66:30:@42804.4]
  assign _T_95268 = _T_95259[8]; // @[OneHot.scala 66:30:@42805.4]
  assign _T_95269 = _T_95259[9]; // @[OneHot.scala 66:30:@42806.4]
  assign _T_95270 = _T_95259[10]; // @[OneHot.scala 66:30:@42807.4]
  assign _T_95271 = _T_95259[11]; // @[OneHot.scala 66:30:@42808.4]
  assign _T_95272 = _T_95259[12]; // @[OneHot.scala 66:30:@42809.4]
  assign _T_95273 = _T_95259[13]; // @[OneHot.scala 66:30:@42810.4]
  assign _T_95274 = _T_95259[14]; // @[OneHot.scala 66:30:@42811.4]
  assign _T_95275 = _T_95259[15]; // @[OneHot.scala 66:30:@42812.4]
  assign _T_95316 = _T_94219 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42830.4]
  assign _T_95317 = _T_94216 ? 16'h4000 : _T_95316; // @[Mux.scala 31:69:@42831.4]
  assign _T_95318 = _T_94213 ? 16'h2000 : _T_95317; // @[Mux.scala 31:69:@42832.4]
  assign _T_95319 = _T_94210 ? 16'h1000 : _T_95318; // @[Mux.scala 31:69:@42833.4]
  assign _T_95320 = _T_94207 ? 16'h800 : _T_95319; // @[Mux.scala 31:69:@42834.4]
  assign _T_95321 = _T_94204 ? 16'h400 : _T_95320; // @[Mux.scala 31:69:@42835.4]
  assign _T_95322 = _T_94201 ? 16'h200 : _T_95321; // @[Mux.scala 31:69:@42836.4]
  assign _T_95323 = _T_94198 ? 16'h100 : _T_95322; // @[Mux.scala 31:69:@42837.4]
  assign _T_95324 = _T_94195 ? 16'h80 : _T_95323; // @[Mux.scala 31:69:@42838.4]
  assign _T_95325 = _T_94192 ? 16'h40 : _T_95324; // @[Mux.scala 31:69:@42839.4]
  assign _T_95326 = _T_94189 ? 16'h20 : _T_95325; // @[Mux.scala 31:69:@42840.4]
  assign _T_95327 = _T_94186 ? 16'h10 : _T_95326; // @[Mux.scala 31:69:@42841.4]
  assign _T_95328 = _T_94183 ? 16'h8 : _T_95327; // @[Mux.scala 31:69:@42842.4]
  assign _T_95329 = _T_94180 ? 16'h4 : _T_95328; // @[Mux.scala 31:69:@42843.4]
  assign _T_95330 = _T_94225 ? 16'h2 : _T_95329; // @[Mux.scala 31:69:@42844.4]
  assign _T_95331 = _T_94222 ? 16'h1 : _T_95330; // @[Mux.scala 31:69:@42845.4]
  assign _T_95332 = _T_95331[0]; // @[OneHot.scala 66:30:@42846.4]
  assign _T_95333 = _T_95331[1]; // @[OneHot.scala 66:30:@42847.4]
  assign _T_95334 = _T_95331[2]; // @[OneHot.scala 66:30:@42848.4]
  assign _T_95335 = _T_95331[3]; // @[OneHot.scala 66:30:@42849.4]
  assign _T_95336 = _T_95331[4]; // @[OneHot.scala 66:30:@42850.4]
  assign _T_95337 = _T_95331[5]; // @[OneHot.scala 66:30:@42851.4]
  assign _T_95338 = _T_95331[6]; // @[OneHot.scala 66:30:@42852.4]
  assign _T_95339 = _T_95331[7]; // @[OneHot.scala 66:30:@42853.4]
  assign _T_95340 = _T_95331[8]; // @[OneHot.scala 66:30:@42854.4]
  assign _T_95341 = _T_95331[9]; // @[OneHot.scala 66:30:@42855.4]
  assign _T_95342 = _T_95331[10]; // @[OneHot.scala 66:30:@42856.4]
  assign _T_95343 = _T_95331[11]; // @[OneHot.scala 66:30:@42857.4]
  assign _T_95344 = _T_95331[12]; // @[OneHot.scala 66:30:@42858.4]
  assign _T_95345 = _T_95331[13]; // @[OneHot.scala 66:30:@42859.4]
  assign _T_95346 = _T_95331[14]; // @[OneHot.scala 66:30:@42860.4]
  assign _T_95347 = _T_95331[15]; // @[OneHot.scala 66:30:@42861.4]
  assign _T_95388 = _T_94222 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@42879.4]
  assign _T_95389 = _T_94219 ? 16'h4000 : _T_95388; // @[Mux.scala 31:69:@42880.4]
  assign _T_95390 = _T_94216 ? 16'h2000 : _T_95389; // @[Mux.scala 31:69:@42881.4]
  assign _T_95391 = _T_94213 ? 16'h1000 : _T_95390; // @[Mux.scala 31:69:@42882.4]
  assign _T_95392 = _T_94210 ? 16'h800 : _T_95391; // @[Mux.scala 31:69:@42883.4]
  assign _T_95393 = _T_94207 ? 16'h400 : _T_95392; // @[Mux.scala 31:69:@42884.4]
  assign _T_95394 = _T_94204 ? 16'h200 : _T_95393; // @[Mux.scala 31:69:@42885.4]
  assign _T_95395 = _T_94201 ? 16'h100 : _T_95394; // @[Mux.scala 31:69:@42886.4]
  assign _T_95396 = _T_94198 ? 16'h80 : _T_95395; // @[Mux.scala 31:69:@42887.4]
  assign _T_95397 = _T_94195 ? 16'h40 : _T_95396; // @[Mux.scala 31:69:@42888.4]
  assign _T_95398 = _T_94192 ? 16'h20 : _T_95397; // @[Mux.scala 31:69:@42889.4]
  assign _T_95399 = _T_94189 ? 16'h10 : _T_95398; // @[Mux.scala 31:69:@42890.4]
  assign _T_95400 = _T_94186 ? 16'h8 : _T_95399; // @[Mux.scala 31:69:@42891.4]
  assign _T_95401 = _T_94183 ? 16'h4 : _T_95400; // @[Mux.scala 31:69:@42892.4]
  assign _T_95402 = _T_94180 ? 16'h2 : _T_95401; // @[Mux.scala 31:69:@42893.4]
  assign _T_95403 = _T_94225 ? 16'h1 : _T_95402; // @[Mux.scala 31:69:@42894.4]
  assign _T_95404 = _T_95403[0]; // @[OneHot.scala 66:30:@42895.4]
  assign _T_95405 = _T_95403[1]; // @[OneHot.scala 66:30:@42896.4]
  assign _T_95406 = _T_95403[2]; // @[OneHot.scala 66:30:@42897.4]
  assign _T_95407 = _T_95403[3]; // @[OneHot.scala 66:30:@42898.4]
  assign _T_95408 = _T_95403[4]; // @[OneHot.scala 66:30:@42899.4]
  assign _T_95409 = _T_95403[5]; // @[OneHot.scala 66:30:@42900.4]
  assign _T_95410 = _T_95403[6]; // @[OneHot.scala 66:30:@42901.4]
  assign _T_95411 = _T_95403[7]; // @[OneHot.scala 66:30:@42902.4]
  assign _T_95412 = _T_95403[8]; // @[OneHot.scala 66:30:@42903.4]
  assign _T_95413 = _T_95403[9]; // @[OneHot.scala 66:30:@42904.4]
  assign _T_95414 = _T_95403[10]; // @[OneHot.scala 66:30:@42905.4]
  assign _T_95415 = _T_95403[11]; // @[OneHot.scala 66:30:@42906.4]
  assign _T_95416 = _T_95403[12]; // @[OneHot.scala 66:30:@42907.4]
  assign _T_95417 = _T_95403[13]; // @[OneHot.scala 66:30:@42908.4]
  assign _T_95418 = _T_95403[14]; // @[OneHot.scala 66:30:@42909.4]
  assign _T_95419 = _T_95403[15]; // @[OneHot.scala 66:30:@42910.4]
  assign _T_95484 = {_T_94331,_T_94330,_T_94329,_T_94328,_T_94327,_T_94326,_T_94325,_T_94324}; // @[Mux.scala 19:72:@42934.4]
  assign _T_95492 = {_T_94339,_T_94338,_T_94337,_T_94336,_T_94335,_T_94334,_T_94333,_T_94332,_T_95484}; // @[Mux.scala 19:72:@42942.4]
  assign _T_95494 = _T_90400 ? _T_95492 : 16'h0; // @[Mux.scala 19:72:@42943.4]
  assign _T_95501 = {_T_94402,_T_94401,_T_94400,_T_94399,_T_94398,_T_94397,_T_94396,_T_94411}; // @[Mux.scala 19:72:@42950.4]
  assign _T_95509 = {_T_94410,_T_94409,_T_94408,_T_94407,_T_94406,_T_94405,_T_94404,_T_94403,_T_95501}; // @[Mux.scala 19:72:@42958.4]
  assign _T_95511 = _T_90401 ? _T_95509 : 16'h0; // @[Mux.scala 19:72:@42959.4]
  assign _T_95518 = {_T_94473,_T_94472,_T_94471,_T_94470,_T_94469,_T_94468,_T_94483,_T_94482}; // @[Mux.scala 19:72:@42966.4]
  assign _T_95526 = {_T_94481,_T_94480,_T_94479,_T_94478,_T_94477,_T_94476,_T_94475,_T_94474,_T_95518}; // @[Mux.scala 19:72:@42974.4]
  assign _T_95528 = _T_90402 ? _T_95526 : 16'h0; // @[Mux.scala 19:72:@42975.4]
  assign _T_95535 = {_T_94544,_T_94543,_T_94542,_T_94541,_T_94540,_T_94555,_T_94554,_T_94553}; // @[Mux.scala 19:72:@42982.4]
  assign _T_95543 = {_T_94552,_T_94551,_T_94550,_T_94549,_T_94548,_T_94547,_T_94546,_T_94545,_T_95535}; // @[Mux.scala 19:72:@42990.4]
  assign _T_95545 = _T_90403 ? _T_95543 : 16'h0; // @[Mux.scala 19:72:@42991.4]
  assign _T_95552 = {_T_94615,_T_94614,_T_94613,_T_94612,_T_94627,_T_94626,_T_94625,_T_94624}; // @[Mux.scala 19:72:@42998.4]
  assign _T_95560 = {_T_94623,_T_94622,_T_94621,_T_94620,_T_94619,_T_94618,_T_94617,_T_94616,_T_95552}; // @[Mux.scala 19:72:@43006.4]
  assign _T_95562 = _T_90404 ? _T_95560 : 16'h0; // @[Mux.scala 19:72:@43007.4]
  assign _T_95569 = {_T_94686,_T_94685,_T_94684,_T_94699,_T_94698,_T_94697,_T_94696,_T_94695}; // @[Mux.scala 19:72:@43014.4]
  assign _T_95577 = {_T_94694,_T_94693,_T_94692,_T_94691,_T_94690,_T_94689,_T_94688,_T_94687,_T_95569}; // @[Mux.scala 19:72:@43022.4]
  assign _T_95579 = _T_90405 ? _T_95577 : 16'h0; // @[Mux.scala 19:72:@43023.4]
  assign _T_95586 = {_T_94757,_T_94756,_T_94771,_T_94770,_T_94769,_T_94768,_T_94767,_T_94766}; // @[Mux.scala 19:72:@43030.4]
  assign _T_95594 = {_T_94765,_T_94764,_T_94763,_T_94762,_T_94761,_T_94760,_T_94759,_T_94758,_T_95586}; // @[Mux.scala 19:72:@43038.4]
  assign _T_95596 = _T_90406 ? _T_95594 : 16'h0; // @[Mux.scala 19:72:@43039.4]
  assign _T_95603 = {_T_94828,_T_94843,_T_94842,_T_94841,_T_94840,_T_94839,_T_94838,_T_94837}; // @[Mux.scala 19:72:@43046.4]
  assign _T_95611 = {_T_94836,_T_94835,_T_94834,_T_94833,_T_94832,_T_94831,_T_94830,_T_94829,_T_95603}; // @[Mux.scala 19:72:@43054.4]
  assign _T_95613 = _T_90407 ? _T_95611 : 16'h0; // @[Mux.scala 19:72:@43055.4]
  assign _T_95620 = {_T_94915,_T_94914,_T_94913,_T_94912,_T_94911,_T_94910,_T_94909,_T_94908}; // @[Mux.scala 19:72:@43062.4]
  assign _T_95628 = {_T_94907,_T_94906,_T_94905,_T_94904,_T_94903,_T_94902,_T_94901,_T_94900,_T_95620}; // @[Mux.scala 19:72:@43070.4]
  assign _T_95630 = _T_90408 ? _T_95628 : 16'h0; // @[Mux.scala 19:72:@43071.4]
  assign _T_95637 = {_T_94986,_T_94985,_T_94984,_T_94983,_T_94982,_T_94981,_T_94980,_T_94979}; // @[Mux.scala 19:72:@43078.4]
  assign _T_95645 = {_T_94978,_T_94977,_T_94976,_T_94975,_T_94974,_T_94973,_T_94972,_T_94987,_T_95637}; // @[Mux.scala 19:72:@43086.4]
  assign _T_95647 = _T_90409 ? _T_95645 : 16'h0; // @[Mux.scala 19:72:@43087.4]
  assign _T_95654 = {_T_95057,_T_95056,_T_95055,_T_95054,_T_95053,_T_95052,_T_95051,_T_95050}; // @[Mux.scala 19:72:@43094.4]
  assign _T_95662 = {_T_95049,_T_95048,_T_95047,_T_95046,_T_95045,_T_95044,_T_95059,_T_95058,_T_95654}; // @[Mux.scala 19:72:@43102.4]
  assign _T_95664 = _T_90410 ? _T_95662 : 16'h0; // @[Mux.scala 19:72:@43103.4]
  assign _T_95671 = {_T_95128,_T_95127,_T_95126,_T_95125,_T_95124,_T_95123,_T_95122,_T_95121}; // @[Mux.scala 19:72:@43110.4]
  assign _T_95679 = {_T_95120,_T_95119,_T_95118,_T_95117,_T_95116,_T_95131,_T_95130,_T_95129,_T_95671}; // @[Mux.scala 19:72:@43118.4]
  assign _T_95681 = _T_90411 ? _T_95679 : 16'h0; // @[Mux.scala 19:72:@43119.4]
  assign _T_95688 = {_T_95199,_T_95198,_T_95197,_T_95196,_T_95195,_T_95194,_T_95193,_T_95192}; // @[Mux.scala 19:72:@43126.4]
  assign _T_95696 = {_T_95191,_T_95190,_T_95189,_T_95188,_T_95203,_T_95202,_T_95201,_T_95200,_T_95688}; // @[Mux.scala 19:72:@43134.4]
  assign _T_95698 = _T_90412 ? _T_95696 : 16'h0; // @[Mux.scala 19:72:@43135.4]
  assign _T_95705 = {_T_95270,_T_95269,_T_95268,_T_95267,_T_95266,_T_95265,_T_95264,_T_95263}; // @[Mux.scala 19:72:@43142.4]
  assign _T_95713 = {_T_95262,_T_95261,_T_95260,_T_95275,_T_95274,_T_95273,_T_95272,_T_95271,_T_95705}; // @[Mux.scala 19:72:@43150.4]
  assign _T_95715 = _T_90413 ? _T_95713 : 16'h0; // @[Mux.scala 19:72:@43151.4]
  assign _T_95722 = {_T_95341,_T_95340,_T_95339,_T_95338,_T_95337,_T_95336,_T_95335,_T_95334}; // @[Mux.scala 19:72:@43158.4]
  assign _T_95730 = {_T_95333,_T_95332,_T_95347,_T_95346,_T_95345,_T_95344,_T_95343,_T_95342,_T_95722}; // @[Mux.scala 19:72:@43166.4]
  assign _T_95732 = _T_90414 ? _T_95730 : 16'h0; // @[Mux.scala 19:72:@43167.4]
  assign _T_95739 = {_T_95412,_T_95411,_T_95410,_T_95409,_T_95408,_T_95407,_T_95406,_T_95405}; // @[Mux.scala 19:72:@43174.4]
  assign _T_95747 = {_T_95404,_T_95419,_T_95418,_T_95417,_T_95416,_T_95415,_T_95414,_T_95413,_T_95739}; // @[Mux.scala 19:72:@43182.4]
  assign _T_95749 = _T_90415 ? _T_95747 : 16'h0; // @[Mux.scala 19:72:@43183.4]
  assign _T_95750 = _T_95494 | _T_95511; // @[Mux.scala 19:72:@43184.4]
  assign _T_95751 = _T_95750 | _T_95528; // @[Mux.scala 19:72:@43185.4]
  assign _T_95752 = _T_95751 | _T_95545; // @[Mux.scala 19:72:@43186.4]
  assign _T_95753 = _T_95752 | _T_95562; // @[Mux.scala 19:72:@43187.4]
  assign _T_95754 = _T_95753 | _T_95579; // @[Mux.scala 19:72:@43188.4]
  assign _T_95755 = _T_95754 | _T_95596; // @[Mux.scala 19:72:@43189.4]
  assign _T_95756 = _T_95755 | _T_95613; // @[Mux.scala 19:72:@43190.4]
  assign _T_95757 = _T_95756 | _T_95630; // @[Mux.scala 19:72:@43191.4]
  assign _T_95758 = _T_95757 | _T_95647; // @[Mux.scala 19:72:@43192.4]
  assign _T_95759 = _T_95758 | _T_95664; // @[Mux.scala 19:72:@43193.4]
  assign _T_95760 = _T_95759 | _T_95681; // @[Mux.scala 19:72:@43194.4]
  assign _T_95761 = _T_95760 | _T_95698; // @[Mux.scala 19:72:@43195.4]
  assign _T_95762 = _T_95761 | _T_95715; // @[Mux.scala 19:72:@43196.4]
  assign _T_95763 = _T_95762 | _T_95732; // @[Mux.scala 19:72:@43197.4]
  assign _T_95764 = _T_95763 | _T_95749; // @[Mux.scala 19:72:@43198.4]
  assign inputPriorityPorts_0_0 = _T_95764[0]; // @[Mux.scala 19:72:@43202.4]
  assign inputPriorityPorts_0_1 = _T_95764[1]; // @[Mux.scala 19:72:@43204.4]
  assign inputPriorityPorts_0_2 = _T_95764[2]; // @[Mux.scala 19:72:@43206.4]
  assign inputPriorityPorts_0_3 = _T_95764[3]; // @[Mux.scala 19:72:@43208.4]
  assign inputPriorityPorts_0_4 = _T_95764[4]; // @[Mux.scala 19:72:@43210.4]
  assign inputPriorityPorts_0_5 = _T_95764[5]; // @[Mux.scala 19:72:@43212.4]
  assign inputPriorityPorts_0_6 = _T_95764[6]; // @[Mux.scala 19:72:@43214.4]
  assign inputPriorityPorts_0_7 = _T_95764[7]; // @[Mux.scala 19:72:@43216.4]
  assign inputPriorityPorts_0_8 = _T_95764[8]; // @[Mux.scala 19:72:@43218.4]
  assign inputPriorityPorts_0_9 = _T_95764[9]; // @[Mux.scala 19:72:@43220.4]
  assign inputPriorityPorts_0_10 = _T_95764[10]; // @[Mux.scala 19:72:@43222.4]
  assign inputPriorityPorts_0_11 = _T_95764[11]; // @[Mux.scala 19:72:@43224.4]
  assign inputPriorityPorts_0_12 = _T_95764[12]; // @[Mux.scala 19:72:@43226.4]
  assign inputPriorityPorts_0_13 = _T_95764[13]; // @[Mux.scala 19:72:@43228.4]
  assign inputPriorityPorts_0_14 = _T_95764[14]; // @[Mux.scala 19:72:@43230.4]
  assign inputPriorityPorts_0_15 = _T_95764[15]; // @[Mux.scala 19:72:@43232.4]
  assign _T_95966 = entriesPorts_0_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43286.4]
  assign _T_95967 = entriesPorts_0_14 ? 16'h4000 : _T_95966; // @[Mux.scala 31:69:@43287.4]
  assign _T_95968 = entriesPorts_0_13 ? 16'h2000 : _T_95967; // @[Mux.scala 31:69:@43288.4]
  assign _T_95969 = entriesPorts_0_12 ? 16'h1000 : _T_95968; // @[Mux.scala 31:69:@43289.4]
  assign _T_95970 = entriesPorts_0_11 ? 16'h800 : _T_95969; // @[Mux.scala 31:69:@43290.4]
  assign _T_95971 = entriesPorts_0_10 ? 16'h400 : _T_95970; // @[Mux.scala 31:69:@43291.4]
  assign _T_95972 = entriesPorts_0_9 ? 16'h200 : _T_95971; // @[Mux.scala 31:69:@43292.4]
  assign _T_95973 = entriesPorts_0_8 ? 16'h100 : _T_95972; // @[Mux.scala 31:69:@43293.4]
  assign _T_95974 = entriesPorts_0_7 ? 16'h80 : _T_95973; // @[Mux.scala 31:69:@43294.4]
  assign _T_95975 = entriesPorts_0_6 ? 16'h40 : _T_95974; // @[Mux.scala 31:69:@43295.4]
  assign _T_95976 = entriesPorts_0_5 ? 16'h20 : _T_95975; // @[Mux.scala 31:69:@43296.4]
  assign _T_95977 = entriesPorts_0_4 ? 16'h10 : _T_95976; // @[Mux.scala 31:69:@43297.4]
  assign _T_95978 = entriesPorts_0_3 ? 16'h8 : _T_95977; // @[Mux.scala 31:69:@43298.4]
  assign _T_95979 = entriesPorts_0_2 ? 16'h4 : _T_95978; // @[Mux.scala 31:69:@43299.4]
  assign _T_95980 = entriesPorts_0_1 ? 16'h2 : _T_95979; // @[Mux.scala 31:69:@43300.4]
  assign _T_95981 = entriesPorts_0_0 ? 16'h1 : _T_95980; // @[Mux.scala 31:69:@43301.4]
  assign _T_95982 = _T_95981[0]; // @[OneHot.scala 66:30:@43302.4]
  assign _T_95983 = _T_95981[1]; // @[OneHot.scala 66:30:@43303.4]
  assign _T_95984 = _T_95981[2]; // @[OneHot.scala 66:30:@43304.4]
  assign _T_95985 = _T_95981[3]; // @[OneHot.scala 66:30:@43305.4]
  assign _T_95986 = _T_95981[4]; // @[OneHot.scala 66:30:@43306.4]
  assign _T_95987 = _T_95981[5]; // @[OneHot.scala 66:30:@43307.4]
  assign _T_95988 = _T_95981[6]; // @[OneHot.scala 66:30:@43308.4]
  assign _T_95989 = _T_95981[7]; // @[OneHot.scala 66:30:@43309.4]
  assign _T_95990 = _T_95981[8]; // @[OneHot.scala 66:30:@43310.4]
  assign _T_95991 = _T_95981[9]; // @[OneHot.scala 66:30:@43311.4]
  assign _T_95992 = _T_95981[10]; // @[OneHot.scala 66:30:@43312.4]
  assign _T_95993 = _T_95981[11]; // @[OneHot.scala 66:30:@43313.4]
  assign _T_95994 = _T_95981[12]; // @[OneHot.scala 66:30:@43314.4]
  assign _T_95995 = _T_95981[13]; // @[OneHot.scala 66:30:@43315.4]
  assign _T_95996 = _T_95981[14]; // @[OneHot.scala 66:30:@43316.4]
  assign _T_95997 = _T_95981[15]; // @[OneHot.scala 66:30:@43317.4]
  assign _T_96038 = entriesPorts_0_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43335.4]
  assign _T_96039 = entriesPorts_0_15 ? 16'h4000 : _T_96038; // @[Mux.scala 31:69:@43336.4]
  assign _T_96040 = entriesPorts_0_14 ? 16'h2000 : _T_96039; // @[Mux.scala 31:69:@43337.4]
  assign _T_96041 = entriesPorts_0_13 ? 16'h1000 : _T_96040; // @[Mux.scala 31:69:@43338.4]
  assign _T_96042 = entriesPorts_0_12 ? 16'h800 : _T_96041; // @[Mux.scala 31:69:@43339.4]
  assign _T_96043 = entriesPorts_0_11 ? 16'h400 : _T_96042; // @[Mux.scala 31:69:@43340.4]
  assign _T_96044 = entriesPorts_0_10 ? 16'h200 : _T_96043; // @[Mux.scala 31:69:@43341.4]
  assign _T_96045 = entriesPorts_0_9 ? 16'h100 : _T_96044; // @[Mux.scala 31:69:@43342.4]
  assign _T_96046 = entriesPorts_0_8 ? 16'h80 : _T_96045; // @[Mux.scala 31:69:@43343.4]
  assign _T_96047 = entriesPorts_0_7 ? 16'h40 : _T_96046; // @[Mux.scala 31:69:@43344.4]
  assign _T_96048 = entriesPorts_0_6 ? 16'h20 : _T_96047; // @[Mux.scala 31:69:@43345.4]
  assign _T_96049 = entriesPorts_0_5 ? 16'h10 : _T_96048; // @[Mux.scala 31:69:@43346.4]
  assign _T_96050 = entriesPorts_0_4 ? 16'h8 : _T_96049; // @[Mux.scala 31:69:@43347.4]
  assign _T_96051 = entriesPorts_0_3 ? 16'h4 : _T_96050; // @[Mux.scala 31:69:@43348.4]
  assign _T_96052 = entriesPorts_0_2 ? 16'h2 : _T_96051; // @[Mux.scala 31:69:@43349.4]
  assign _T_96053 = entriesPorts_0_1 ? 16'h1 : _T_96052; // @[Mux.scala 31:69:@43350.4]
  assign _T_96054 = _T_96053[0]; // @[OneHot.scala 66:30:@43351.4]
  assign _T_96055 = _T_96053[1]; // @[OneHot.scala 66:30:@43352.4]
  assign _T_96056 = _T_96053[2]; // @[OneHot.scala 66:30:@43353.4]
  assign _T_96057 = _T_96053[3]; // @[OneHot.scala 66:30:@43354.4]
  assign _T_96058 = _T_96053[4]; // @[OneHot.scala 66:30:@43355.4]
  assign _T_96059 = _T_96053[5]; // @[OneHot.scala 66:30:@43356.4]
  assign _T_96060 = _T_96053[6]; // @[OneHot.scala 66:30:@43357.4]
  assign _T_96061 = _T_96053[7]; // @[OneHot.scala 66:30:@43358.4]
  assign _T_96062 = _T_96053[8]; // @[OneHot.scala 66:30:@43359.4]
  assign _T_96063 = _T_96053[9]; // @[OneHot.scala 66:30:@43360.4]
  assign _T_96064 = _T_96053[10]; // @[OneHot.scala 66:30:@43361.4]
  assign _T_96065 = _T_96053[11]; // @[OneHot.scala 66:30:@43362.4]
  assign _T_96066 = _T_96053[12]; // @[OneHot.scala 66:30:@43363.4]
  assign _T_96067 = _T_96053[13]; // @[OneHot.scala 66:30:@43364.4]
  assign _T_96068 = _T_96053[14]; // @[OneHot.scala 66:30:@43365.4]
  assign _T_96069 = _T_96053[15]; // @[OneHot.scala 66:30:@43366.4]
  assign _T_96110 = entriesPorts_0_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43384.4]
  assign _T_96111 = entriesPorts_0_0 ? 16'h4000 : _T_96110; // @[Mux.scala 31:69:@43385.4]
  assign _T_96112 = entriesPorts_0_15 ? 16'h2000 : _T_96111; // @[Mux.scala 31:69:@43386.4]
  assign _T_96113 = entriesPorts_0_14 ? 16'h1000 : _T_96112; // @[Mux.scala 31:69:@43387.4]
  assign _T_96114 = entriesPorts_0_13 ? 16'h800 : _T_96113; // @[Mux.scala 31:69:@43388.4]
  assign _T_96115 = entriesPorts_0_12 ? 16'h400 : _T_96114; // @[Mux.scala 31:69:@43389.4]
  assign _T_96116 = entriesPorts_0_11 ? 16'h200 : _T_96115; // @[Mux.scala 31:69:@43390.4]
  assign _T_96117 = entriesPorts_0_10 ? 16'h100 : _T_96116; // @[Mux.scala 31:69:@43391.4]
  assign _T_96118 = entriesPorts_0_9 ? 16'h80 : _T_96117; // @[Mux.scala 31:69:@43392.4]
  assign _T_96119 = entriesPorts_0_8 ? 16'h40 : _T_96118; // @[Mux.scala 31:69:@43393.4]
  assign _T_96120 = entriesPorts_0_7 ? 16'h20 : _T_96119; // @[Mux.scala 31:69:@43394.4]
  assign _T_96121 = entriesPorts_0_6 ? 16'h10 : _T_96120; // @[Mux.scala 31:69:@43395.4]
  assign _T_96122 = entriesPorts_0_5 ? 16'h8 : _T_96121; // @[Mux.scala 31:69:@43396.4]
  assign _T_96123 = entriesPorts_0_4 ? 16'h4 : _T_96122; // @[Mux.scala 31:69:@43397.4]
  assign _T_96124 = entriesPorts_0_3 ? 16'h2 : _T_96123; // @[Mux.scala 31:69:@43398.4]
  assign _T_96125 = entriesPorts_0_2 ? 16'h1 : _T_96124; // @[Mux.scala 31:69:@43399.4]
  assign _T_96126 = _T_96125[0]; // @[OneHot.scala 66:30:@43400.4]
  assign _T_96127 = _T_96125[1]; // @[OneHot.scala 66:30:@43401.4]
  assign _T_96128 = _T_96125[2]; // @[OneHot.scala 66:30:@43402.4]
  assign _T_96129 = _T_96125[3]; // @[OneHot.scala 66:30:@43403.4]
  assign _T_96130 = _T_96125[4]; // @[OneHot.scala 66:30:@43404.4]
  assign _T_96131 = _T_96125[5]; // @[OneHot.scala 66:30:@43405.4]
  assign _T_96132 = _T_96125[6]; // @[OneHot.scala 66:30:@43406.4]
  assign _T_96133 = _T_96125[7]; // @[OneHot.scala 66:30:@43407.4]
  assign _T_96134 = _T_96125[8]; // @[OneHot.scala 66:30:@43408.4]
  assign _T_96135 = _T_96125[9]; // @[OneHot.scala 66:30:@43409.4]
  assign _T_96136 = _T_96125[10]; // @[OneHot.scala 66:30:@43410.4]
  assign _T_96137 = _T_96125[11]; // @[OneHot.scala 66:30:@43411.4]
  assign _T_96138 = _T_96125[12]; // @[OneHot.scala 66:30:@43412.4]
  assign _T_96139 = _T_96125[13]; // @[OneHot.scala 66:30:@43413.4]
  assign _T_96140 = _T_96125[14]; // @[OneHot.scala 66:30:@43414.4]
  assign _T_96141 = _T_96125[15]; // @[OneHot.scala 66:30:@43415.4]
  assign _T_96182 = entriesPorts_0_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43433.4]
  assign _T_96183 = entriesPorts_0_1 ? 16'h4000 : _T_96182; // @[Mux.scala 31:69:@43434.4]
  assign _T_96184 = entriesPorts_0_0 ? 16'h2000 : _T_96183; // @[Mux.scala 31:69:@43435.4]
  assign _T_96185 = entriesPorts_0_15 ? 16'h1000 : _T_96184; // @[Mux.scala 31:69:@43436.4]
  assign _T_96186 = entriesPorts_0_14 ? 16'h800 : _T_96185; // @[Mux.scala 31:69:@43437.4]
  assign _T_96187 = entriesPorts_0_13 ? 16'h400 : _T_96186; // @[Mux.scala 31:69:@43438.4]
  assign _T_96188 = entriesPorts_0_12 ? 16'h200 : _T_96187; // @[Mux.scala 31:69:@43439.4]
  assign _T_96189 = entriesPorts_0_11 ? 16'h100 : _T_96188; // @[Mux.scala 31:69:@43440.4]
  assign _T_96190 = entriesPorts_0_10 ? 16'h80 : _T_96189; // @[Mux.scala 31:69:@43441.4]
  assign _T_96191 = entriesPorts_0_9 ? 16'h40 : _T_96190; // @[Mux.scala 31:69:@43442.4]
  assign _T_96192 = entriesPorts_0_8 ? 16'h20 : _T_96191; // @[Mux.scala 31:69:@43443.4]
  assign _T_96193 = entriesPorts_0_7 ? 16'h10 : _T_96192; // @[Mux.scala 31:69:@43444.4]
  assign _T_96194 = entriesPorts_0_6 ? 16'h8 : _T_96193; // @[Mux.scala 31:69:@43445.4]
  assign _T_96195 = entriesPorts_0_5 ? 16'h4 : _T_96194; // @[Mux.scala 31:69:@43446.4]
  assign _T_96196 = entriesPorts_0_4 ? 16'h2 : _T_96195; // @[Mux.scala 31:69:@43447.4]
  assign _T_96197 = entriesPorts_0_3 ? 16'h1 : _T_96196; // @[Mux.scala 31:69:@43448.4]
  assign _T_96198 = _T_96197[0]; // @[OneHot.scala 66:30:@43449.4]
  assign _T_96199 = _T_96197[1]; // @[OneHot.scala 66:30:@43450.4]
  assign _T_96200 = _T_96197[2]; // @[OneHot.scala 66:30:@43451.4]
  assign _T_96201 = _T_96197[3]; // @[OneHot.scala 66:30:@43452.4]
  assign _T_96202 = _T_96197[4]; // @[OneHot.scala 66:30:@43453.4]
  assign _T_96203 = _T_96197[5]; // @[OneHot.scala 66:30:@43454.4]
  assign _T_96204 = _T_96197[6]; // @[OneHot.scala 66:30:@43455.4]
  assign _T_96205 = _T_96197[7]; // @[OneHot.scala 66:30:@43456.4]
  assign _T_96206 = _T_96197[8]; // @[OneHot.scala 66:30:@43457.4]
  assign _T_96207 = _T_96197[9]; // @[OneHot.scala 66:30:@43458.4]
  assign _T_96208 = _T_96197[10]; // @[OneHot.scala 66:30:@43459.4]
  assign _T_96209 = _T_96197[11]; // @[OneHot.scala 66:30:@43460.4]
  assign _T_96210 = _T_96197[12]; // @[OneHot.scala 66:30:@43461.4]
  assign _T_96211 = _T_96197[13]; // @[OneHot.scala 66:30:@43462.4]
  assign _T_96212 = _T_96197[14]; // @[OneHot.scala 66:30:@43463.4]
  assign _T_96213 = _T_96197[15]; // @[OneHot.scala 66:30:@43464.4]
  assign _T_96254 = entriesPorts_0_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43482.4]
  assign _T_96255 = entriesPorts_0_2 ? 16'h4000 : _T_96254; // @[Mux.scala 31:69:@43483.4]
  assign _T_96256 = entriesPorts_0_1 ? 16'h2000 : _T_96255; // @[Mux.scala 31:69:@43484.4]
  assign _T_96257 = entriesPorts_0_0 ? 16'h1000 : _T_96256; // @[Mux.scala 31:69:@43485.4]
  assign _T_96258 = entriesPorts_0_15 ? 16'h800 : _T_96257; // @[Mux.scala 31:69:@43486.4]
  assign _T_96259 = entriesPorts_0_14 ? 16'h400 : _T_96258; // @[Mux.scala 31:69:@43487.4]
  assign _T_96260 = entriesPorts_0_13 ? 16'h200 : _T_96259; // @[Mux.scala 31:69:@43488.4]
  assign _T_96261 = entriesPorts_0_12 ? 16'h100 : _T_96260; // @[Mux.scala 31:69:@43489.4]
  assign _T_96262 = entriesPorts_0_11 ? 16'h80 : _T_96261; // @[Mux.scala 31:69:@43490.4]
  assign _T_96263 = entriesPorts_0_10 ? 16'h40 : _T_96262; // @[Mux.scala 31:69:@43491.4]
  assign _T_96264 = entriesPorts_0_9 ? 16'h20 : _T_96263; // @[Mux.scala 31:69:@43492.4]
  assign _T_96265 = entriesPorts_0_8 ? 16'h10 : _T_96264; // @[Mux.scala 31:69:@43493.4]
  assign _T_96266 = entriesPorts_0_7 ? 16'h8 : _T_96265; // @[Mux.scala 31:69:@43494.4]
  assign _T_96267 = entriesPorts_0_6 ? 16'h4 : _T_96266; // @[Mux.scala 31:69:@43495.4]
  assign _T_96268 = entriesPorts_0_5 ? 16'h2 : _T_96267; // @[Mux.scala 31:69:@43496.4]
  assign _T_96269 = entriesPorts_0_4 ? 16'h1 : _T_96268; // @[Mux.scala 31:69:@43497.4]
  assign _T_96270 = _T_96269[0]; // @[OneHot.scala 66:30:@43498.4]
  assign _T_96271 = _T_96269[1]; // @[OneHot.scala 66:30:@43499.4]
  assign _T_96272 = _T_96269[2]; // @[OneHot.scala 66:30:@43500.4]
  assign _T_96273 = _T_96269[3]; // @[OneHot.scala 66:30:@43501.4]
  assign _T_96274 = _T_96269[4]; // @[OneHot.scala 66:30:@43502.4]
  assign _T_96275 = _T_96269[5]; // @[OneHot.scala 66:30:@43503.4]
  assign _T_96276 = _T_96269[6]; // @[OneHot.scala 66:30:@43504.4]
  assign _T_96277 = _T_96269[7]; // @[OneHot.scala 66:30:@43505.4]
  assign _T_96278 = _T_96269[8]; // @[OneHot.scala 66:30:@43506.4]
  assign _T_96279 = _T_96269[9]; // @[OneHot.scala 66:30:@43507.4]
  assign _T_96280 = _T_96269[10]; // @[OneHot.scala 66:30:@43508.4]
  assign _T_96281 = _T_96269[11]; // @[OneHot.scala 66:30:@43509.4]
  assign _T_96282 = _T_96269[12]; // @[OneHot.scala 66:30:@43510.4]
  assign _T_96283 = _T_96269[13]; // @[OneHot.scala 66:30:@43511.4]
  assign _T_96284 = _T_96269[14]; // @[OneHot.scala 66:30:@43512.4]
  assign _T_96285 = _T_96269[15]; // @[OneHot.scala 66:30:@43513.4]
  assign _T_96326 = entriesPorts_0_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43531.4]
  assign _T_96327 = entriesPorts_0_3 ? 16'h4000 : _T_96326; // @[Mux.scala 31:69:@43532.4]
  assign _T_96328 = entriesPorts_0_2 ? 16'h2000 : _T_96327; // @[Mux.scala 31:69:@43533.4]
  assign _T_96329 = entriesPorts_0_1 ? 16'h1000 : _T_96328; // @[Mux.scala 31:69:@43534.4]
  assign _T_96330 = entriesPorts_0_0 ? 16'h800 : _T_96329; // @[Mux.scala 31:69:@43535.4]
  assign _T_96331 = entriesPorts_0_15 ? 16'h400 : _T_96330; // @[Mux.scala 31:69:@43536.4]
  assign _T_96332 = entriesPorts_0_14 ? 16'h200 : _T_96331; // @[Mux.scala 31:69:@43537.4]
  assign _T_96333 = entriesPorts_0_13 ? 16'h100 : _T_96332; // @[Mux.scala 31:69:@43538.4]
  assign _T_96334 = entriesPorts_0_12 ? 16'h80 : _T_96333; // @[Mux.scala 31:69:@43539.4]
  assign _T_96335 = entriesPorts_0_11 ? 16'h40 : _T_96334; // @[Mux.scala 31:69:@43540.4]
  assign _T_96336 = entriesPorts_0_10 ? 16'h20 : _T_96335; // @[Mux.scala 31:69:@43541.4]
  assign _T_96337 = entriesPorts_0_9 ? 16'h10 : _T_96336; // @[Mux.scala 31:69:@43542.4]
  assign _T_96338 = entriesPorts_0_8 ? 16'h8 : _T_96337; // @[Mux.scala 31:69:@43543.4]
  assign _T_96339 = entriesPorts_0_7 ? 16'h4 : _T_96338; // @[Mux.scala 31:69:@43544.4]
  assign _T_96340 = entriesPorts_0_6 ? 16'h2 : _T_96339; // @[Mux.scala 31:69:@43545.4]
  assign _T_96341 = entriesPorts_0_5 ? 16'h1 : _T_96340; // @[Mux.scala 31:69:@43546.4]
  assign _T_96342 = _T_96341[0]; // @[OneHot.scala 66:30:@43547.4]
  assign _T_96343 = _T_96341[1]; // @[OneHot.scala 66:30:@43548.4]
  assign _T_96344 = _T_96341[2]; // @[OneHot.scala 66:30:@43549.4]
  assign _T_96345 = _T_96341[3]; // @[OneHot.scala 66:30:@43550.4]
  assign _T_96346 = _T_96341[4]; // @[OneHot.scala 66:30:@43551.4]
  assign _T_96347 = _T_96341[5]; // @[OneHot.scala 66:30:@43552.4]
  assign _T_96348 = _T_96341[6]; // @[OneHot.scala 66:30:@43553.4]
  assign _T_96349 = _T_96341[7]; // @[OneHot.scala 66:30:@43554.4]
  assign _T_96350 = _T_96341[8]; // @[OneHot.scala 66:30:@43555.4]
  assign _T_96351 = _T_96341[9]; // @[OneHot.scala 66:30:@43556.4]
  assign _T_96352 = _T_96341[10]; // @[OneHot.scala 66:30:@43557.4]
  assign _T_96353 = _T_96341[11]; // @[OneHot.scala 66:30:@43558.4]
  assign _T_96354 = _T_96341[12]; // @[OneHot.scala 66:30:@43559.4]
  assign _T_96355 = _T_96341[13]; // @[OneHot.scala 66:30:@43560.4]
  assign _T_96356 = _T_96341[14]; // @[OneHot.scala 66:30:@43561.4]
  assign _T_96357 = _T_96341[15]; // @[OneHot.scala 66:30:@43562.4]
  assign _T_96398 = entriesPorts_0_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43580.4]
  assign _T_96399 = entriesPorts_0_4 ? 16'h4000 : _T_96398; // @[Mux.scala 31:69:@43581.4]
  assign _T_96400 = entriesPorts_0_3 ? 16'h2000 : _T_96399; // @[Mux.scala 31:69:@43582.4]
  assign _T_96401 = entriesPorts_0_2 ? 16'h1000 : _T_96400; // @[Mux.scala 31:69:@43583.4]
  assign _T_96402 = entriesPorts_0_1 ? 16'h800 : _T_96401; // @[Mux.scala 31:69:@43584.4]
  assign _T_96403 = entriesPorts_0_0 ? 16'h400 : _T_96402; // @[Mux.scala 31:69:@43585.4]
  assign _T_96404 = entriesPorts_0_15 ? 16'h200 : _T_96403; // @[Mux.scala 31:69:@43586.4]
  assign _T_96405 = entriesPorts_0_14 ? 16'h100 : _T_96404; // @[Mux.scala 31:69:@43587.4]
  assign _T_96406 = entriesPorts_0_13 ? 16'h80 : _T_96405; // @[Mux.scala 31:69:@43588.4]
  assign _T_96407 = entriesPorts_0_12 ? 16'h40 : _T_96406; // @[Mux.scala 31:69:@43589.4]
  assign _T_96408 = entriesPorts_0_11 ? 16'h20 : _T_96407; // @[Mux.scala 31:69:@43590.4]
  assign _T_96409 = entriesPorts_0_10 ? 16'h10 : _T_96408; // @[Mux.scala 31:69:@43591.4]
  assign _T_96410 = entriesPorts_0_9 ? 16'h8 : _T_96409; // @[Mux.scala 31:69:@43592.4]
  assign _T_96411 = entriesPorts_0_8 ? 16'h4 : _T_96410; // @[Mux.scala 31:69:@43593.4]
  assign _T_96412 = entriesPorts_0_7 ? 16'h2 : _T_96411; // @[Mux.scala 31:69:@43594.4]
  assign _T_96413 = entriesPorts_0_6 ? 16'h1 : _T_96412; // @[Mux.scala 31:69:@43595.4]
  assign _T_96414 = _T_96413[0]; // @[OneHot.scala 66:30:@43596.4]
  assign _T_96415 = _T_96413[1]; // @[OneHot.scala 66:30:@43597.4]
  assign _T_96416 = _T_96413[2]; // @[OneHot.scala 66:30:@43598.4]
  assign _T_96417 = _T_96413[3]; // @[OneHot.scala 66:30:@43599.4]
  assign _T_96418 = _T_96413[4]; // @[OneHot.scala 66:30:@43600.4]
  assign _T_96419 = _T_96413[5]; // @[OneHot.scala 66:30:@43601.4]
  assign _T_96420 = _T_96413[6]; // @[OneHot.scala 66:30:@43602.4]
  assign _T_96421 = _T_96413[7]; // @[OneHot.scala 66:30:@43603.4]
  assign _T_96422 = _T_96413[8]; // @[OneHot.scala 66:30:@43604.4]
  assign _T_96423 = _T_96413[9]; // @[OneHot.scala 66:30:@43605.4]
  assign _T_96424 = _T_96413[10]; // @[OneHot.scala 66:30:@43606.4]
  assign _T_96425 = _T_96413[11]; // @[OneHot.scala 66:30:@43607.4]
  assign _T_96426 = _T_96413[12]; // @[OneHot.scala 66:30:@43608.4]
  assign _T_96427 = _T_96413[13]; // @[OneHot.scala 66:30:@43609.4]
  assign _T_96428 = _T_96413[14]; // @[OneHot.scala 66:30:@43610.4]
  assign _T_96429 = _T_96413[15]; // @[OneHot.scala 66:30:@43611.4]
  assign _T_96470 = entriesPorts_0_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43629.4]
  assign _T_96471 = entriesPorts_0_5 ? 16'h4000 : _T_96470; // @[Mux.scala 31:69:@43630.4]
  assign _T_96472 = entriesPorts_0_4 ? 16'h2000 : _T_96471; // @[Mux.scala 31:69:@43631.4]
  assign _T_96473 = entriesPorts_0_3 ? 16'h1000 : _T_96472; // @[Mux.scala 31:69:@43632.4]
  assign _T_96474 = entriesPorts_0_2 ? 16'h800 : _T_96473; // @[Mux.scala 31:69:@43633.4]
  assign _T_96475 = entriesPorts_0_1 ? 16'h400 : _T_96474; // @[Mux.scala 31:69:@43634.4]
  assign _T_96476 = entriesPorts_0_0 ? 16'h200 : _T_96475; // @[Mux.scala 31:69:@43635.4]
  assign _T_96477 = entriesPorts_0_15 ? 16'h100 : _T_96476; // @[Mux.scala 31:69:@43636.4]
  assign _T_96478 = entriesPorts_0_14 ? 16'h80 : _T_96477; // @[Mux.scala 31:69:@43637.4]
  assign _T_96479 = entriesPorts_0_13 ? 16'h40 : _T_96478; // @[Mux.scala 31:69:@43638.4]
  assign _T_96480 = entriesPorts_0_12 ? 16'h20 : _T_96479; // @[Mux.scala 31:69:@43639.4]
  assign _T_96481 = entriesPorts_0_11 ? 16'h10 : _T_96480; // @[Mux.scala 31:69:@43640.4]
  assign _T_96482 = entriesPorts_0_10 ? 16'h8 : _T_96481; // @[Mux.scala 31:69:@43641.4]
  assign _T_96483 = entriesPorts_0_9 ? 16'h4 : _T_96482; // @[Mux.scala 31:69:@43642.4]
  assign _T_96484 = entriesPorts_0_8 ? 16'h2 : _T_96483; // @[Mux.scala 31:69:@43643.4]
  assign _T_96485 = entriesPorts_0_7 ? 16'h1 : _T_96484; // @[Mux.scala 31:69:@43644.4]
  assign _T_96486 = _T_96485[0]; // @[OneHot.scala 66:30:@43645.4]
  assign _T_96487 = _T_96485[1]; // @[OneHot.scala 66:30:@43646.4]
  assign _T_96488 = _T_96485[2]; // @[OneHot.scala 66:30:@43647.4]
  assign _T_96489 = _T_96485[3]; // @[OneHot.scala 66:30:@43648.4]
  assign _T_96490 = _T_96485[4]; // @[OneHot.scala 66:30:@43649.4]
  assign _T_96491 = _T_96485[5]; // @[OneHot.scala 66:30:@43650.4]
  assign _T_96492 = _T_96485[6]; // @[OneHot.scala 66:30:@43651.4]
  assign _T_96493 = _T_96485[7]; // @[OneHot.scala 66:30:@43652.4]
  assign _T_96494 = _T_96485[8]; // @[OneHot.scala 66:30:@43653.4]
  assign _T_96495 = _T_96485[9]; // @[OneHot.scala 66:30:@43654.4]
  assign _T_96496 = _T_96485[10]; // @[OneHot.scala 66:30:@43655.4]
  assign _T_96497 = _T_96485[11]; // @[OneHot.scala 66:30:@43656.4]
  assign _T_96498 = _T_96485[12]; // @[OneHot.scala 66:30:@43657.4]
  assign _T_96499 = _T_96485[13]; // @[OneHot.scala 66:30:@43658.4]
  assign _T_96500 = _T_96485[14]; // @[OneHot.scala 66:30:@43659.4]
  assign _T_96501 = _T_96485[15]; // @[OneHot.scala 66:30:@43660.4]
  assign _T_96542 = entriesPorts_0_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43678.4]
  assign _T_96543 = entriesPorts_0_6 ? 16'h4000 : _T_96542; // @[Mux.scala 31:69:@43679.4]
  assign _T_96544 = entriesPorts_0_5 ? 16'h2000 : _T_96543; // @[Mux.scala 31:69:@43680.4]
  assign _T_96545 = entriesPorts_0_4 ? 16'h1000 : _T_96544; // @[Mux.scala 31:69:@43681.4]
  assign _T_96546 = entriesPorts_0_3 ? 16'h800 : _T_96545; // @[Mux.scala 31:69:@43682.4]
  assign _T_96547 = entriesPorts_0_2 ? 16'h400 : _T_96546; // @[Mux.scala 31:69:@43683.4]
  assign _T_96548 = entriesPorts_0_1 ? 16'h200 : _T_96547; // @[Mux.scala 31:69:@43684.4]
  assign _T_96549 = entriesPorts_0_0 ? 16'h100 : _T_96548; // @[Mux.scala 31:69:@43685.4]
  assign _T_96550 = entriesPorts_0_15 ? 16'h80 : _T_96549; // @[Mux.scala 31:69:@43686.4]
  assign _T_96551 = entriesPorts_0_14 ? 16'h40 : _T_96550; // @[Mux.scala 31:69:@43687.4]
  assign _T_96552 = entriesPorts_0_13 ? 16'h20 : _T_96551; // @[Mux.scala 31:69:@43688.4]
  assign _T_96553 = entriesPorts_0_12 ? 16'h10 : _T_96552; // @[Mux.scala 31:69:@43689.4]
  assign _T_96554 = entriesPorts_0_11 ? 16'h8 : _T_96553; // @[Mux.scala 31:69:@43690.4]
  assign _T_96555 = entriesPorts_0_10 ? 16'h4 : _T_96554; // @[Mux.scala 31:69:@43691.4]
  assign _T_96556 = entriesPorts_0_9 ? 16'h2 : _T_96555; // @[Mux.scala 31:69:@43692.4]
  assign _T_96557 = entriesPorts_0_8 ? 16'h1 : _T_96556; // @[Mux.scala 31:69:@43693.4]
  assign _T_96558 = _T_96557[0]; // @[OneHot.scala 66:30:@43694.4]
  assign _T_96559 = _T_96557[1]; // @[OneHot.scala 66:30:@43695.4]
  assign _T_96560 = _T_96557[2]; // @[OneHot.scala 66:30:@43696.4]
  assign _T_96561 = _T_96557[3]; // @[OneHot.scala 66:30:@43697.4]
  assign _T_96562 = _T_96557[4]; // @[OneHot.scala 66:30:@43698.4]
  assign _T_96563 = _T_96557[5]; // @[OneHot.scala 66:30:@43699.4]
  assign _T_96564 = _T_96557[6]; // @[OneHot.scala 66:30:@43700.4]
  assign _T_96565 = _T_96557[7]; // @[OneHot.scala 66:30:@43701.4]
  assign _T_96566 = _T_96557[8]; // @[OneHot.scala 66:30:@43702.4]
  assign _T_96567 = _T_96557[9]; // @[OneHot.scala 66:30:@43703.4]
  assign _T_96568 = _T_96557[10]; // @[OneHot.scala 66:30:@43704.4]
  assign _T_96569 = _T_96557[11]; // @[OneHot.scala 66:30:@43705.4]
  assign _T_96570 = _T_96557[12]; // @[OneHot.scala 66:30:@43706.4]
  assign _T_96571 = _T_96557[13]; // @[OneHot.scala 66:30:@43707.4]
  assign _T_96572 = _T_96557[14]; // @[OneHot.scala 66:30:@43708.4]
  assign _T_96573 = _T_96557[15]; // @[OneHot.scala 66:30:@43709.4]
  assign _T_96614 = entriesPorts_0_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43727.4]
  assign _T_96615 = entriesPorts_0_7 ? 16'h4000 : _T_96614; // @[Mux.scala 31:69:@43728.4]
  assign _T_96616 = entriesPorts_0_6 ? 16'h2000 : _T_96615; // @[Mux.scala 31:69:@43729.4]
  assign _T_96617 = entriesPorts_0_5 ? 16'h1000 : _T_96616; // @[Mux.scala 31:69:@43730.4]
  assign _T_96618 = entriesPorts_0_4 ? 16'h800 : _T_96617; // @[Mux.scala 31:69:@43731.4]
  assign _T_96619 = entriesPorts_0_3 ? 16'h400 : _T_96618; // @[Mux.scala 31:69:@43732.4]
  assign _T_96620 = entriesPorts_0_2 ? 16'h200 : _T_96619; // @[Mux.scala 31:69:@43733.4]
  assign _T_96621 = entriesPorts_0_1 ? 16'h100 : _T_96620; // @[Mux.scala 31:69:@43734.4]
  assign _T_96622 = entriesPorts_0_0 ? 16'h80 : _T_96621; // @[Mux.scala 31:69:@43735.4]
  assign _T_96623 = entriesPorts_0_15 ? 16'h40 : _T_96622; // @[Mux.scala 31:69:@43736.4]
  assign _T_96624 = entriesPorts_0_14 ? 16'h20 : _T_96623; // @[Mux.scala 31:69:@43737.4]
  assign _T_96625 = entriesPorts_0_13 ? 16'h10 : _T_96624; // @[Mux.scala 31:69:@43738.4]
  assign _T_96626 = entriesPorts_0_12 ? 16'h8 : _T_96625; // @[Mux.scala 31:69:@43739.4]
  assign _T_96627 = entriesPorts_0_11 ? 16'h4 : _T_96626; // @[Mux.scala 31:69:@43740.4]
  assign _T_96628 = entriesPorts_0_10 ? 16'h2 : _T_96627; // @[Mux.scala 31:69:@43741.4]
  assign _T_96629 = entriesPorts_0_9 ? 16'h1 : _T_96628; // @[Mux.scala 31:69:@43742.4]
  assign _T_96630 = _T_96629[0]; // @[OneHot.scala 66:30:@43743.4]
  assign _T_96631 = _T_96629[1]; // @[OneHot.scala 66:30:@43744.4]
  assign _T_96632 = _T_96629[2]; // @[OneHot.scala 66:30:@43745.4]
  assign _T_96633 = _T_96629[3]; // @[OneHot.scala 66:30:@43746.4]
  assign _T_96634 = _T_96629[4]; // @[OneHot.scala 66:30:@43747.4]
  assign _T_96635 = _T_96629[5]; // @[OneHot.scala 66:30:@43748.4]
  assign _T_96636 = _T_96629[6]; // @[OneHot.scala 66:30:@43749.4]
  assign _T_96637 = _T_96629[7]; // @[OneHot.scala 66:30:@43750.4]
  assign _T_96638 = _T_96629[8]; // @[OneHot.scala 66:30:@43751.4]
  assign _T_96639 = _T_96629[9]; // @[OneHot.scala 66:30:@43752.4]
  assign _T_96640 = _T_96629[10]; // @[OneHot.scala 66:30:@43753.4]
  assign _T_96641 = _T_96629[11]; // @[OneHot.scala 66:30:@43754.4]
  assign _T_96642 = _T_96629[12]; // @[OneHot.scala 66:30:@43755.4]
  assign _T_96643 = _T_96629[13]; // @[OneHot.scala 66:30:@43756.4]
  assign _T_96644 = _T_96629[14]; // @[OneHot.scala 66:30:@43757.4]
  assign _T_96645 = _T_96629[15]; // @[OneHot.scala 66:30:@43758.4]
  assign _T_96686 = entriesPorts_0_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43776.4]
  assign _T_96687 = entriesPorts_0_8 ? 16'h4000 : _T_96686; // @[Mux.scala 31:69:@43777.4]
  assign _T_96688 = entriesPorts_0_7 ? 16'h2000 : _T_96687; // @[Mux.scala 31:69:@43778.4]
  assign _T_96689 = entriesPorts_0_6 ? 16'h1000 : _T_96688; // @[Mux.scala 31:69:@43779.4]
  assign _T_96690 = entriesPorts_0_5 ? 16'h800 : _T_96689; // @[Mux.scala 31:69:@43780.4]
  assign _T_96691 = entriesPorts_0_4 ? 16'h400 : _T_96690; // @[Mux.scala 31:69:@43781.4]
  assign _T_96692 = entriesPorts_0_3 ? 16'h200 : _T_96691; // @[Mux.scala 31:69:@43782.4]
  assign _T_96693 = entriesPorts_0_2 ? 16'h100 : _T_96692; // @[Mux.scala 31:69:@43783.4]
  assign _T_96694 = entriesPorts_0_1 ? 16'h80 : _T_96693; // @[Mux.scala 31:69:@43784.4]
  assign _T_96695 = entriesPorts_0_0 ? 16'h40 : _T_96694; // @[Mux.scala 31:69:@43785.4]
  assign _T_96696 = entriesPorts_0_15 ? 16'h20 : _T_96695; // @[Mux.scala 31:69:@43786.4]
  assign _T_96697 = entriesPorts_0_14 ? 16'h10 : _T_96696; // @[Mux.scala 31:69:@43787.4]
  assign _T_96698 = entriesPorts_0_13 ? 16'h8 : _T_96697; // @[Mux.scala 31:69:@43788.4]
  assign _T_96699 = entriesPorts_0_12 ? 16'h4 : _T_96698; // @[Mux.scala 31:69:@43789.4]
  assign _T_96700 = entriesPorts_0_11 ? 16'h2 : _T_96699; // @[Mux.scala 31:69:@43790.4]
  assign _T_96701 = entriesPorts_0_10 ? 16'h1 : _T_96700; // @[Mux.scala 31:69:@43791.4]
  assign _T_96702 = _T_96701[0]; // @[OneHot.scala 66:30:@43792.4]
  assign _T_96703 = _T_96701[1]; // @[OneHot.scala 66:30:@43793.4]
  assign _T_96704 = _T_96701[2]; // @[OneHot.scala 66:30:@43794.4]
  assign _T_96705 = _T_96701[3]; // @[OneHot.scala 66:30:@43795.4]
  assign _T_96706 = _T_96701[4]; // @[OneHot.scala 66:30:@43796.4]
  assign _T_96707 = _T_96701[5]; // @[OneHot.scala 66:30:@43797.4]
  assign _T_96708 = _T_96701[6]; // @[OneHot.scala 66:30:@43798.4]
  assign _T_96709 = _T_96701[7]; // @[OneHot.scala 66:30:@43799.4]
  assign _T_96710 = _T_96701[8]; // @[OneHot.scala 66:30:@43800.4]
  assign _T_96711 = _T_96701[9]; // @[OneHot.scala 66:30:@43801.4]
  assign _T_96712 = _T_96701[10]; // @[OneHot.scala 66:30:@43802.4]
  assign _T_96713 = _T_96701[11]; // @[OneHot.scala 66:30:@43803.4]
  assign _T_96714 = _T_96701[12]; // @[OneHot.scala 66:30:@43804.4]
  assign _T_96715 = _T_96701[13]; // @[OneHot.scala 66:30:@43805.4]
  assign _T_96716 = _T_96701[14]; // @[OneHot.scala 66:30:@43806.4]
  assign _T_96717 = _T_96701[15]; // @[OneHot.scala 66:30:@43807.4]
  assign _T_96758 = entriesPorts_0_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43825.4]
  assign _T_96759 = entriesPorts_0_9 ? 16'h4000 : _T_96758; // @[Mux.scala 31:69:@43826.4]
  assign _T_96760 = entriesPorts_0_8 ? 16'h2000 : _T_96759; // @[Mux.scala 31:69:@43827.4]
  assign _T_96761 = entriesPorts_0_7 ? 16'h1000 : _T_96760; // @[Mux.scala 31:69:@43828.4]
  assign _T_96762 = entriesPorts_0_6 ? 16'h800 : _T_96761; // @[Mux.scala 31:69:@43829.4]
  assign _T_96763 = entriesPorts_0_5 ? 16'h400 : _T_96762; // @[Mux.scala 31:69:@43830.4]
  assign _T_96764 = entriesPorts_0_4 ? 16'h200 : _T_96763; // @[Mux.scala 31:69:@43831.4]
  assign _T_96765 = entriesPorts_0_3 ? 16'h100 : _T_96764; // @[Mux.scala 31:69:@43832.4]
  assign _T_96766 = entriesPorts_0_2 ? 16'h80 : _T_96765; // @[Mux.scala 31:69:@43833.4]
  assign _T_96767 = entriesPorts_0_1 ? 16'h40 : _T_96766; // @[Mux.scala 31:69:@43834.4]
  assign _T_96768 = entriesPorts_0_0 ? 16'h20 : _T_96767; // @[Mux.scala 31:69:@43835.4]
  assign _T_96769 = entriesPorts_0_15 ? 16'h10 : _T_96768; // @[Mux.scala 31:69:@43836.4]
  assign _T_96770 = entriesPorts_0_14 ? 16'h8 : _T_96769; // @[Mux.scala 31:69:@43837.4]
  assign _T_96771 = entriesPorts_0_13 ? 16'h4 : _T_96770; // @[Mux.scala 31:69:@43838.4]
  assign _T_96772 = entriesPorts_0_12 ? 16'h2 : _T_96771; // @[Mux.scala 31:69:@43839.4]
  assign _T_96773 = entriesPorts_0_11 ? 16'h1 : _T_96772; // @[Mux.scala 31:69:@43840.4]
  assign _T_96774 = _T_96773[0]; // @[OneHot.scala 66:30:@43841.4]
  assign _T_96775 = _T_96773[1]; // @[OneHot.scala 66:30:@43842.4]
  assign _T_96776 = _T_96773[2]; // @[OneHot.scala 66:30:@43843.4]
  assign _T_96777 = _T_96773[3]; // @[OneHot.scala 66:30:@43844.4]
  assign _T_96778 = _T_96773[4]; // @[OneHot.scala 66:30:@43845.4]
  assign _T_96779 = _T_96773[5]; // @[OneHot.scala 66:30:@43846.4]
  assign _T_96780 = _T_96773[6]; // @[OneHot.scala 66:30:@43847.4]
  assign _T_96781 = _T_96773[7]; // @[OneHot.scala 66:30:@43848.4]
  assign _T_96782 = _T_96773[8]; // @[OneHot.scala 66:30:@43849.4]
  assign _T_96783 = _T_96773[9]; // @[OneHot.scala 66:30:@43850.4]
  assign _T_96784 = _T_96773[10]; // @[OneHot.scala 66:30:@43851.4]
  assign _T_96785 = _T_96773[11]; // @[OneHot.scala 66:30:@43852.4]
  assign _T_96786 = _T_96773[12]; // @[OneHot.scala 66:30:@43853.4]
  assign _T_96787 = _T_96773[13]; // @[OneHot.scala 66:30:@43854.4]
  assign _T_96788 = _T_96773[14]; // @[OneHot.scala 66:30:@43855.4]
  assign _T_96789 = _T_96773[15]; // @[OneHot.scala 66:30:@43856.4]
  assign _T_96830 = entriesPorts_0_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43874.4]
  assign _T_96831 = entriesPorts_0_10 ? 16'h4000 : _T_96830; // @[Mux.scala 31:69:@43875.4]
  assign _T_96832 = entriesPorts_0_9 ? 16'h2000 : _T_96831; // @[Mux.scala 31:69:@43876.4]
  assign _T_96833 = entriesPorts_0_8 ? 16'h1000 : _T_96832; // @[Mux.scala 31:69:@43877.4]
  assign _T_96834 = entriesPorts_0_7 ? 16'h800 : _T_96833; // @[Mux.scala 31:69:@43878.4]
  assign _T_96835 = entriesPorts_0_6 ? 16'h400 : _T_96834; // @[Mux.scala 31:69:@43879.4]
  assign _T_96836 = entriesPorts_0_5 ? 16'h200 : _T_96835; // @[Mux.scala 31:69:@43880.4]
  assign _T_96837 = entriesPorts_0_4 ? 16'h100 : _T_96836; // @[Mux.scala 31:69:@43881.4]
  assign _T_96838 = entriesPorts_0_3 ? 16'h80 : _T_96837; // @[Mux.scala 31:69:@43882.4]
  assign _T_96839 = entriesPorts_0_2 ? 16'h40 : _T_96838; // @[Mux.scala 31:69:@43883.4]
  assign _T_96840 = entriesPorts_0_1 ? 16'h20 : _T_96839; // @[Mux.scala 31:69:@43884.4]
  assign _T_96841 = entriesPorts_0_0 ? 16'h10 : _T_96840; // @[Mux.scala 31:69:@43885.4]
  assign _T_96842 = entriesPorts_0_15 ? 16'h8 : _T_96841; // @[Mux.scala 31:69:@43886.4]
  assign _T_96843 = entriesPorts_0_14 ? 16'h4 : _T_96842; // @[Mux.scala 31:69:@43887.4]
  assign _T_96844 = entriesPorts_0_13 ? 16'h2 : _T_96843; // @[Mux.scala 31:69:@43888.4]
  assign _T_96845 = entriesPorts_0_12 ? 16'h1 : _T_96844; // @[Mux.scala 31:69:@43889.4]
  assign _T_96846 = _T_96845[0]; // @[OneHot.scala 66:30:@43890.4]
  assign _T_96847 = _T_96845[1]; // @[OneHot.scala 66:30:@43891.4]
  assign _T_96848 = _T_96845[2]; // @[OneHot.scala 66:30:@43892.4]
  assign _T_96849 = _T_96845[3]; // @[OneHot.scala 66:30:@43893.4]
  assign _T_96850 = _T_96845[4]; // @[OneHot.scala 66:30:@43894.4]
  assign _T_96851 = _T_96845[5]; // @[OneHot.scala 66:30:@43895.4]
  assign _T_96852 = _T_96845[6]; // @[OneHot.scala 66:30:@43896.4]
  assign _T_96853 = _T_96845[7]; // @[OneHot.scala 66:30:@43897.4]
  assign _T_96854 = _T_96845[8]; // @[OneHot.scala 66:30:@43898.4]
  assign _T_96855 = _T_96845[9]; // @[OneHot.scala 66:30:@43899.4]
  assign _T_96856 = _T_96845[10]; // @[OneHot.scala 66:30:@43900.4]
  assign _T_96857 = _T_96845[11]; // @[OneHot.scala 66:30:@43901.4]
  assign _T_96858 = _T_96845[12]; // @[OneHot.scala 66:30:@43902.4]
  assign _T_96859 = _T_96845[13]; // @[OneHot.scala 66:30:@43903.4]
  assign _T_96860 = _T_96845[14]; // @[OneHot.scala 66:30:@43904.4]
  assign _T_96861 = _T_96845[15]; // @[OneHot.scala 66:30:@43905.4]
  assign _T_96902 = entriesPorts_0_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43923.4]
  assign _T_96903 = entriesPorts_0_11 ? 16'h4000 : _T_96902; // @[Mux.scala 31:69:@43924.4]
  assign _T_96904 = entriesPorts_0_10 ? 16'h2000 : _T_96903; // @[Mux.scala 31:69:@43925.4]
  assign _T_96905 = entriesPorts_0_9 ? 16'h1000 : _T_96904; // @[Mux.scala 31:69:@43926.4]
  assign _T_96906 = entriesPorts_0_8 ? 16'h800 : _T_96905; // @[Mux.scala 31:69:@43927.4]
  assign _T_96907 = entriesPorts_0_7 ? 16'h400 : _T_96906; // @[Mux.scala 31:69:@43928.4]
  assign _T_96908 = entriesPorts_0_6 ? 16'h200 : _T_96907; // @[Mux.scala 31:69:@43929.4]
  assign _T_96909 = entriesPorts_0_5 ? 16'h100 : _T_96908; // @[Mux.scala 31:69:@43930.4]
  assign _T_96910 = entriesPorts_0_4 ? 16'h80 : _T_96909; // @[Mux.scala 31:69:@43931.4]
  assign _T_96911 = entriesPorts_0_3 ? 16'h40 : _T_96910; // @[Mux.scala 31:69:@43932.4]
  assign _T_96912 = entriesPorts_0_2 ? 16'h20 : _T_96911; // @[Mux.scala 31:69:@43933.4]
  assign _T_96913 = entriesPorts_0_1 ? 16'h10 : _T_96912; // @[Mux.scala 31:69:@43934.4]
  assign _T_96914 = entriesPorts_0_0 ? 16'h8 : _T_96913; // @[Mux.scala 31:69:@43935.4]
  assign _T_96915 = entriesPorts_0_15 ? 16'h4 : _T_96914; // @[Mux.scala 31:69:@43936.4]
  assign _T_96916 = entriesPorts_0_14 ? 16'h2 : _T_96915; // @[Mux.scala 31:69:@43937.4]
  assign _T_96917 = entriesPorts_0_13 ? 16'h1 : _T_96916; // @[Mux.scala 31:69:@43938.4]
  assign _T_96918 = _T_96917[0]; // @[OneHot.scala 66:30:@43939.4]
  assign _T_96919 = _T_96917[1]; // @[OneHot.scala 66:30:@43940.4]
  assign _T_96920 = _T_96917[2]; // @[OneHot.scala 66:30:@43941.4]
  assign _T_96921 = _T_96917[3]; // @[OneHot.scala 66:30:@43942.4]
  assign _T_96922 = _T_96917[4]; // @[OneHot.scala 66:30:@43943.4]
  assign _T_96923 = _T_96917[5]; // @[OneHot.scala 66:30:@43944.4]
  assign _T_96924 = _T_96917[6]; // @[OneHot.scala 66:30:@43945.4]
  assign _T_96925 = _T_96917[7]; // @[OneHot.scala 66:30:@43946.4]
  assign _T_96926 = _T_96917[8]; // @[OneHot.scala 66:30:@43947.4]
  assign _T_96927 = _T_96917[9]; // @[OneHot.scala 66:30:@43948.4]
  assign _T_96928 = _T_96917[10]; // @[OneHot.scala 66:30:@43949.4]
  assign _T_96929 = _T_96917[11]; // @[OneHot.scala 66:30:@43950.4]
  assign _T_96930 = _T_96917[12]; // @[OneHot.scala 66:30:@43951.4]
  assign _T_96931 = _T_96917[13]; // @[OneHot.scala 66:30:@43952.4]
  assign _T_96932 = _T_96917[14]; // @[OneHot.scala 66:30:@43953.4]
  assign _T_96933 = _T_96917[15]; // @[OneHot.scala 66:30:@43954.4]
  assign _T_96974 = entriesPorts_0_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@43972.4]
  assign _T_96975 = entriesPorts_0_12 ? 16'h4000 : _T_96974; // @[Mux.scala 31:69:@43973.4]
  assign _T_96976 = entriesPorts_0_11 ? 16'h2000 : _T_96975; // @[Mux.scala 31:69:@43974.4]
  assign _T_96977 = entriesPorts_0_10 ? 16'h1000 : _T_96976; // @[Mux.scala 31:69:@43975.4]
  assign _T_96978 = entriesPorts_0_9 ? 16'h800 : _T_96977; // @[Mux.scala 31:69:@43976.4]
  assign _T_96979 = entriesPorts_0_8 ? 16'h400 : _T_96978; // @[Mux.scala 31:69:@43977.4]
  assign _T_96980 = entriesPorts_0_7 ? 16'h200 : _T_96979; // @[Mux.scala 31:69:@43978.4]
  assign _T_96981 = entriesPorts_0_6 ? 16'h100 : _T_96980; // @[Mux.scala 31:69:@43979.4]
  assign _T_96982 = entriesPorts_0_5 ? 16'h80 : _T_96981; // @[Mux.scala 31:69:@43980.4]
  assign _T_96983 = entriesPorts_0_4 ? 16'h40 : _T_96982; // @[Mux.scala 31:69:@43981.4]
  assign _T_96984 = entriesPorts_0_3 ? 16'h20 : _T_96983; // @[Mux.scala 31:69:@43982.4]
  assign _T_96985 = entriesPorts_0_2 ? 16'h10 : _T_96984; // @[Mux.scala 31:69:@43983.4]
  assign _T_96986 = entriesPorts_0_1 ? 16'h8 : _T_96985; // @[Mux.scala 31:69:@43984.4]
  assign _T_96987 = entriesPorts_0_0 ? 16'h4 : _T_96986; // @[Mux.scala 31:69:@43985.4]
  assign _T_96988 = entriesPorts_0_15 ? 16'h2 : _T_96987; // @[Mux.scala 31:69:@43986.4]
  assign _T_96989 = entriesPorts_0_14 ? 16'h1 : _T_96988; // @[Mux.scala 31:69:@43987.4]
  assign _T_96990 = _T_96989[0]; // @[OneHot.scala 66:30:@43988.4]
  assign _T_96991 = _T_96989[1]; // @[OneHot.scala 66:30:@43989.4]
  assign _T_96992 = _T_96989[2]; // @[OneHot.scala 66:30:@43990.4]
  assign _T_96993 = _T_96989[3]; // @[OneHot.scala 66:30:@43991.4]
  assign _T_96994 = _T_96989[4]; // @[OneHot.scala 66:30:@43992.4]
  assign _T_96995 = _T_96989[5]; // @[OneHot.scala 66:30:@43993.4]
  assign _T_96996 = _T_96989[6]; // @[OneHot.scala 66:30:@43994.4]
  assign _T_96997 = _T_96989[7]; // @[OneHot.scala 66:30:@43995.4]
  assign _T_96998 = _T_96989[8]; // @[OneHot.scala 66:30:@43996.4]
  assign _T_96999 = _T_96989[9]; // @[OneHot.scala 66:30:@43997.4]
  assign _T_97000 = _T_96989[10]; // @[OneHot.scala 66:30:@43998.4]
  assign _T_97001 = _T_96989[11]; // @[OneHot.scala 66:30:@43999.4]
  assign _T_97002 = _T_96989[12]; // @[OneHot.scala 66:30:@44000.4]
  assign _T_97003 = _T_96989[13]; // @[OneHot.scala 66:30:@44001.4]
  assign _T_97004 = _T_96989[14]; // @[OneHot.scala 66:30:@44002.4]
  assign _T_97005 = _T_96989[15]; // @[OneHot.scala 66:30:@44003.4]
  assign _T_97046 = entriesPorts_0_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@44021.4]
  assign _T_97047 = entriesPorts_0_13 ? 16'h4000 : _T_97046; // @[Mux.scala 31:69:@44022.4]
  assign _T_97048 = entriesPorts_0_12 ? 16'h2000 : _T_97047; // @[Mux.scala 31:69:@44023.4]
  assign _T_97049 = entriesPorts_0_11 ? 16'h1000 : _T_97048; // @[Mux.scala 31:69:@44024.4]
  assign _T_97050 = entriesPorts_0_10 ? 16'h800 : _T_97049; // @[Mux.scala 31:69:@44025.4]
  assign _T_97051 = entriesPorts_0_9 ? 16'h400 : _T_97050; // @[Mux.scala 31:69:@44026.4]
  assign _T_97052 = entriesPorts_0_8 ? 16'h200 : _T_97051; // @[Mux.scala 31:69:@44027.4]
  assign _T_97053 = entriesPorts_0_7 ? 16'h100 : _T_97052; // @[Mux.scala 31:69:@44028.4]
  assign _T_97054 = entriesPorts_0_6 ? 16'h80 : _T_97053; // @[Mux.scala 31:69:@44029.4]
  assign _T_97055 = entriesPorts_0_5 ? 16'h40 : _T_97054; // @[Mux.scala 31:69:@44030.4]
  assign _T_97056 = entriesPorts_0_4 ? 16'h20 : _T_97055; // @[Mux.scala 31:69:@44031.4]
  assign _T_97057 = entriesPorts_0_3 ? 16'h10 : _T_97056; // @[Mux.scala 31:69:@44032.4]
  assign _T_97058 = entriesPorts_0_2 ? 16'h8 : _T_97057; // @[Mux.scala 31:69:@44033.4]
  assign _T_97059 = entriesPorts_0_1 ? 16'h4 : _T_97058; // @[Mux.scala 31:69:@44034.4]
  assign _T_97060 = entriesPorts_0_0 ? 16'h2 : _T_97059; // @[Mux.scala 31:69:@44035.4]
  assign _T_97061 = entriesPorts_0_15 ? 16'h1 : _T_97060; // @[Mux.scala 31:69:@44036.4]
  assign _T_97062 = _T_97061[0]; // @[OneHot.scala 66:30:@44037.4]
  assign _T_97063 = _T_97061[1]; // @[OneHot.scala 66:30:@44038.4]
  assign _T_97064 = _T_97061[2]; // @[OneHot.scala 66:30:@44039.4]
  assign _T_97065 = _T_97061[3]; // @[OneHot.scala 66:30:@44040.4]
  assign _T_97066 = _T_97061[4]; // @[OneHot.scala 66:30:@44041.4]
  assign _T_97067 = _T_97061[5]; // @[OneHot.scala 66:30:@44042.4]
  assign _T_97068 = _T_97061[6]; // @[OneHot.scala 66:30:@44043.4]
  assign _T_97069 = _T_97061[7]; // @[OneHot.scala 66:30:@44044.4]
  assign _T_97070 = _T_97061[8]; // @[OneHot.scala 66:30:@44045.4]
  assign _T_97071 = _T_97061[9]; // @[OneHot.scala 66:30:@44046.4]
  assign _T_97072 = _T_97061[10]; // @[OneHot.scala 66:30:@44047.4]
  assign _T_97073 = _T_97061[11]; // @[OneHot.scala 66:30:@44048.4]
  assign _T_97074 = _T_97061[12]; // @[OneHot.scala 66:30:@44049.4]
  assign _T_97075 = _T_97061[13]; // @[OneHot.scala 66:30:@44050.4]
  assign _T_97076 = _T_97061[14]; // @[OneHot.scala 66:30:@44051.4]
  assign _T_97077 = _T_97061[15]; // @[OneHot.scala 66:30:@44052.4]
  assign _T_97142 = {_T_95989,_T_95988,_T_95987,_T_95986,_T_95985,_T_95984,_T_95983,_T_95982}; // @[Mux.scala 19:72:@44076.4]
  assign _T_97150 = {_T_95997,_T_95996,_T_95995,_T_95994,_T_95993,_T_95992,_T_95991,_T_95990,_T_97142}; // @[Mux.scala 19:72:@44084.4]
  assign _T_97152 = _T_90400 ? _T_97150 : 16'h0; // @[Mux.scala 19:72:@44085.4]
  assign _T_97159 = {_T_96060,_T_96059,_T_96058,_T_96057,_T_96056,_T_96055,_T_96054,_T_96069}; // @[Mux.scala 19:72:@44092.4]
  assign _T_97167 = {_T_96068,_T_96067,_T_96066,_T_96065,_T_96064,_T_96063,_T_96062,_T_96061,_T_97159}; // @[Mux.scala 19:72:@44100.4]
  assign _T_97169 = _T_90401 ? _T_97167 : 16'h0; // @[Mux.scala 19:72:@44101.4]
  assign _T_97176 = {_T_96131,_T_96130,_T_96129,_T_96128,_T_96127,_T_96126,_T_96141,_T_96140}; // @[Mux.scala 19:72:@44108.4]
  assign _T_97184 = {_T_96139,_T_96138,_T_96137,_T_96136,_T_96135,_T_96134,_T_96133,_T_96132,_T_97176}; // @[Mux.scala 19:72:@44116.4]
  assign _T_97186 = _T_90402 ? _T_97184 : 16'h0; // @[Mux.scala 19:72:@44117.4]
  assign _T_97193 = {_T_96202,_T_96201,_T_96200,_T_96199,_T_96198,_T_96213,_T_96212,_T_96211}; // @[Mux.scala 19:72:@44124.4]
  assign _T_97201 = {_T_96210,_T_96209,_T_96208,_T_96207,_T_96206,_T_96205,_T_96204,_T_96203,_T_97193}; // @[Mux.scala 19:72:@44132.4]
  assign _T_97203 = _T_90403 ? _T_97201 : 16'h0; // @[Mux.scala 19:72:@44133.4]
  assign _T_97210 = {_T_96273,_T_96272,_T_96271,_T_96270,_T_96285,_T_96284,_T_96283,_T_96282}; // @[Mux.scala 19:72:@44140.4]
  assign _T_97218 = {_T_96281,_T_96280,_T_96279,_T_96278,_T_96277,_T_96276,_T_96275,_T_96274,_T_97210}; // @[Mux.scala 19:72:@44148.4]
  assign _T_97220 = _T_90404 ? _T_97218 : 16'h0; // @[Mux.scala 19:72:@44149.4]
  assign _T_97227 = {_T_96344,_T_96343,_T_96342,_T_96357,_T_96356,_T_96355,_T_96354,_T_96353}; // @[Mux.scala 19:72:@44156.4]
  assign _T_97235 = {_T_96352,_T_96351,_T_96350,_T_96349,_T_96348,_T_96347,_T_96346,_T_96345,_T_97227}; // @[Mux.scala 19:72:@44164.4]
  assign _T_97237 = _T_90405 ? _T_97235 : 16'h0; // @[Mux.scala 19:72:@44165.4]
  assign _T_97244 = {_T_96415,_T_96414,_T_96429,_T_96428,_T_96427,_T_96426,_T_96425,_T_96424}; // @[Mux.scala 19:72:@44172.4]
  assign _T_97252 = {_T_96423,_T_96422,_T_96421,_T_96420,_T_96419,_T_96418,_T_96417,_T_96416,_T_97244}; // @[Mux.scala 19:72:@44180.4]
  assign _T_97254 = _T_90406 ? _T_97252 : 16'h0; // @[Mux.scala 19:72:@44181.4]
  assign _T_97261 = {_T_96486,_T_96501,_T_96500,_T_96499,_T_96498,_T_96497,_T_96496,_T_96495}; // @[Mux.scala 19:72:@44188.4]
  assign _T_97269 = {_T_96494,_T_96493,_T_96492,_T_96491,_T_96490,_T_96489,_T_96488,_T_96487,_T_97261}; // @[Mux.scala 19:72:@44196.4]
  assign _T_97271 = _T_90407 ? _T_97269 : 16'h0; // @[Mux.scala 19:72:@44197.4]
  assign _T_97278 = {_T_96573,_T_96572,_T_96571,_T_96570,_T_96569,_T_96568,_T_96567,_T_96566}; // @[Mux.scala 19:72:@44204.4]
  assign _T_97286 = {_T_96565,_T_96564,_T_96563,_T_96562,_T_96561,_T_96560,_T_96559,_T_96558,_T_97278}; // @[Mux.scala 19:72:@44212.4]
  assign _T_97288 = _T_90408 ? _T_97286 : 16'h0; // @[Mux.scala 19:72:@44213.4]
  assign _T_97295 = {_T_96644,_T_96643,_T_96642,_T_96641,_T_96640,_T_96639,_T_96638,_T_96637}; // @[Mux.scala 19:72:@44220.4]
  assign _T_97303 = {_T_96636,_T_96635,_T_96634,_T_96633,_T_96632,_T_96631,_T_96630,_T_96645,_T_97295}; // @[Mux.scala 19:72:@44228.4]
  assign _T_97305 = _T_90409 ? _T_97303 : 16'h0; // @[Mux.scala 19:72:@44229.4]
  assign _T_97312 = {_T_96715,_T_96714,_T_96713,_T_96712,_T_96711,_T_96710,_T_96709,_T_96708}; // @[Mux.scala 19:72:@44236.4]
  assign _T_97320 = {_T_96707,_T_96706,_T_96705,_T_96704,_T_96703,_T_96702,_T_96717,_T_96716,_T_97312}; // @[Mux.scala 19:72:@44244.4]
  assign _T_97322 = _T_90410 ? _T_97320 : 16'h0; // @[Mux.scala 19:72:@44245.4]
  assign _T_97329 = {_T_96786,_T_96785,_T_96784,_T_96783,_T_96782,_T_96781,_T_96780,_T_96779}; // @[Mux.scala 19:72:@44252.4]
  assign _T_97337 = {_T_96778,_T_96777,_T_96776,_T_96775,_T_96774,_T_96789,_T_96788,_T_96787,_T_97329}; // @[Mux.scala 19:72:@44260.4]
  assign _T_97339 = _T_90411 ? _T_97337 : 16'h0; // @[Mux.scala 19:72:@44261.4]
  assign _T_97346 = {_T_96857,_T_96856,_T_96855,_T_96854,_T_96853,_T_96852,_T_96851,_T_96850}; // @[Mux.scala 19:72:@44268.4]
  assign _T_97354 = {_T_96849,_T_96848,_T_96847,_T_96846,_T_96861,_T_96860,_T_96859,_T_96858,_T_97346}; // @[Mux.scala 19:72:@44276.4]
  assign _T_97356 = _T_90412 ? _T_97354 : 16'h0; // @[Mux.scala 19:72:@44277.4]
  assign _T_97363 = {_T_96928,_T_96927,_T_96926,_T_96925,_T_96924,_T_96923,_T_96922,_T_96921}; // @[Mux.scala 19:72:@44284.4]
  assign _T_97371 = {_T_96920,_T_96919,_T_96918,_T_96933,_T_96932,_T_96931,_T_96930,_T_96929,_T_97363}; // @[Mux.scala 19:72:@44292.4]
  assign _T_97373 = _T_90413 ? _T_97371 : 16'h0; // @[Mux.scala 19:72:@44293.4]
  assign _T_97380 = {_T_96999,_T_96998,_T_96997,_T_96996,_T_96995,_T_96994,_T_96993,_T_96992}; // @[Mux.scala 19:72:@44300.4]
  assign _T_97388 = {_T_96991,_T_96990,_T_97005,_T_97004,_T_97003,_T_97002,_T_97001,_T_97000,_T_97380}; // @[Mux.scala 19:72:@44308.4]
  assign _T_97390 = _T_90414 ? _T_97388 : 16'h0; // @[Mux.scala 19:72:@44309.4]
  assign _T_97397 = {_T_97070,_T_97069,_T_97068,_T_97067,_T_97066,_T_97065,_T_97064,_T_97063}; // @[Mux.scala 19:72:@44316.4]
  assign _T_97405 = {_T_97062,_T_97077,_T_97076,_T_97075,_T_97074,_T_97073,_T_97072,_T_97071,_T_97397}; // @[Mux.scala 19:72:@44324.4]
  assign _T_97407 = _T_90415 ? _T_97405 : 16'h0; // @[Mux.scala 19:72:@44325.4]
  assign _T_97408 = _T_97152 | _T_97169; // @[Mux.scala 19:72:@44326.4]
  assign _T_97409 = _T_97408 | _T_97186; // @[Mux.scala 19:72:@44327.4]
  assign _T_97410 = _T_97409 | _T_97203; // @[Mux.scala 19:72:@44328.4]
  assign _T_97411 = _T_97410 | _T_97220; // @[Mux.scala 19:72:@44329.4]
  assign _T_97412 = _T_97411 | _T_97237; // @[Mux.scala 19:72:@44330.4]
  assign _T_97413 = _T_97412 | _T_97254; // @[Mux.scala 19:72:@44331.4]
  assign _T_97414 = _T_97413 | _T_97271; // @[Mux.scala 19:72:@44332.4]
  assign _T_97415 = _T_97414 | _T_97288; // @[Mux.scala 19:72:@44333.4]
  assign _T_97416 = _T_97415 | _T_97305; // @[Mux.scala 19:72:@44334.4]
  assign _T_97417 = _T_97416 | _T_97322; // @[Mux.scala 19:72:@44335.4]
  assign _T_97418 = _T_97417 | _T_97339; // @[Mux.scala 19:72:@44336.4]
  assign _T_97419 = _T_97418 | _T_97356; // @[Mux.scala 19:72:@44337.4]
  assign _T_97420 = _T_97419 | _T_97373; // @[Mux.scala 19:72:@44338.4]
  assign _T_97421 = _T_97420 | _T_97390; // @[Mux.scala 19:72:@44339.4]
  assign _T_97422 = _T_97421 | _T_97407; // @[Mux.scala 19:72:@44340.4]
  assign outputPriorityPorts_0_0 = _T_97422[0]; // @[Mux.scala 19:72:@44344.4]
  assign outputPriorityPorts_0_1 = _T_97422[1]; // @[Mux.scala 19:72:@44346.4]
  assign outputPriorityPorts_0_2 = _T_97422[2]; // @[Mux.scala 19:72:@44348.4]
  assign outputPriorityPorts_0_3 = _T_97422[3]; // @[Mux.scala 19:72:@44350.4]
  assign outputPriorityPorts_0_4 = _T_97422[4]; // @[Mux.scala 19:72:@44352.4]
  assign outputPriorityPorts_0_5 = _T_97422[5]; // @[Mux.scala 19:72:@44354.4]
  assign outputPriorityPorts_0_6 = _T_97422[6]; // @[Mux.scala 19:72:@44356.4]
  assign outputPriorityPorts_0_7 = _T_97422[7]; // @[Mux.scala 19:72:@44358.4]
  assign outputPriorityPorts_0_8 = _T_97422[8]; // @[Mux.scala 19:72:@44360.4]
  assign outputPriorityPorts_0_9 = _T_97422[9]; // @[Mux.scala 19:72:@44362.4]
  assign outputPriorityPorts_0_10 = _T_97422[10]; // @[Mux.scala 19:72:@44364.4]
  assign outputPriorityPorts_0_11 = _T_97422[11]; // @[Mux.scala 19:72:@44366.4]
  assign outputPriorityPorts_0_12 = _T_97422[12]; // @[Mux.scala 19:72:@44368.4]
  assign outputPriorityPorts_0_13 = _T_97422[13]; // @[Mux.scala 19:72:@44370.4]
  assign outputPriorityPorts_0_14 = _T_97422[14]; // @[Mux.scala 19:72:@44372.4]
  assign outputPriorityPorts_0_15 = _T_97422[15]; // @[Mux.scala 19:72:@44374.4]
  assign _T_97565 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44396.6]
  assign _GEN_2114 = _T_97565 ? io_addrFromLoadPorts_0 : addrQ_0; // @[LoadQueue.scala 314:36:@44400.6]
  assign _GEN_2115 = _T_97565 ? 1'h1 : addrKnown_0; // @[LoadQueue.scala 314:36:@44400.6]
  assign _GEN_2116 = initBits_0 ? 1'h0 : _GEN_2115; // @[LoadQueue.scala 308:34:@44392.4]
  assign _GEN_2117 = initBits_0 ? addrQ_0 : _GEN_2114; // @[LoadQueue.scala 308:34:@44392.4]
  assign _T_97580 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44409.6]
  assign _GEN_2118 = _T_97580 ? io_addrFromLoadPorts_0 : addrQ_1; // @[LoadQueue.scala 314:36:@44413.6]
  assign _GEN_2119 = _T_97580 ? 1'h1 : addrKnown_1; // @[LoadQueue.scala 314:36:@44413.6]
  assign _GEN_2120 = initBits_1 ? 1'h0 : _GEN_2119; // @[LoadQueue.scala 308:34:@44405.4]
  assign _GEN_2121 = initBits_1 ? addrQ_1 : _GEN_2118; // @[LoadQueue.scala 308:34:@44405.4]
  assign _T_97595 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44422.6]
  assign _GEN_2122 = _T_97595 ? io_addrFromLoadPorts_0 : addrQ_2; // @[LoadQueue.scala 314:36:@44426.6]
  assign _GEN_2123 = _T_97595 ? 1'h1 : addrKnown_2; // @[LoadQueue.scala 314:36:@44426.6]
  assign _GEN_2124 = initBits_2 ? 1'h0 : _GEN_2123; // @[LoadQueue.scala 308:34:@44418.4]
  assign _GEN_2125 = initBits_2 ? addrQ_2 : _GEN_2122; // @[LoadQueue.scala 308:34:@44418.4]
  assign _T_97610 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44435.6]
  assign _GEN_2126 = _T_97610 ? io_addrFromLoadPorts_0 : addrQ_3; // @[LoadQueue.scala 314:36:@44439.6]
  assign _GEN_2127 = _T_97610 ? 1'h1 : addrKnown_3; // @[LoadQueue.scala 314:36:@44439.6]
  assign _GEN_2128 = initBits_3 ? 1'h0 : _GEN_2127; // @[LoadQueue.scala 308:34:@44431.4]
  assign _GEN_2129 = initBits_3 ? addrQ_3 : _GEN_2126; // @[LoadQueue.scala 308:34:@44431.4]
  assign _T_97625 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44448.6]
  assign _GEN_2130 = _T_97625 ? io_addrFromLoadPorts_0 : addrQ_4; // @[LoadQueue.scala 314:36:@44452.6]
  assign _GEN_2131 = _T_97625 ? 1'h1 : addrKnown_4; // @[LoadQueue.scala 314:36:@44452.6]
  assign _GEN_2132 = initBits_4 ? 1'h0 : _GEN_2131; // @[LoadQueue.scala 308:34:@44444.4]
  assign _GEN_2133 = initBits_4 ? addrQ_4 : _GEN_2130; // @[LoadQueue.scala 308:34:@44444.4]
  assign _T_97640 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44461.6]
  assign _GEN_2134 = _T_97640 ? io_addrFromLoadPorts_0 : addrQ_5; // @[LoadQueue.scala 314:36:@44465.6]
  assign _GEN_2135 = _T_97640 ? 1'h1 : addrKnown_5; // @[LoadQueue.scala 314:36:@44465.6]
  assign _GEN_2136 = initBits_5 ? 1'h0 : _GEN_2135; // @[LoadQueue.scala 308:34:@44457.4]
  assign _GEN_2137 = initBits_5 ? addrQ_5 : _GEN_2134; // @[LoadQueue.scala 308:34:@44457.4]
  assign _T_97655 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44474.6]
  assign _GEN_2138 = _T_97655 ? io_addrFromLoadPorts_0 : addrQ_6; // @[LoadQueue.scala 314:36:@44478.6]
  assign _GEN_2139 = _T_97655 ? 1'h1 : addrKnown_6; // @[LoadQueue.scala 314:36:@44478.6]
  assign _GEN_2140 = initBits_6 ? 1'h0 : _GEN_2139; // @[LoadQueue.scala 308:34:@44470.4]
  assign _GEN_2141 = initBits_6 ? addrQ_6 : _GEN_2138; // @[LoadQueue.scala 308:34:@44470.4]
  assign _T_97670 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44487.6]
  assign _GEN_2142 = _T_97670 ? io_addrFromLoadPorts_0 : addrQ_7; // @[LoadQueue.scala 314:36:@44491.6]
  assign _GEN_2143 = _T_97670 ? 1'h1 : addrKnown_7; // @[LoadQueue.scala 314:36:@44491.6]
  assign _GEN_2144 = initBits_7 ? 1'h0 : _GEN_2143; // @[LoadQueue.scala 308:34:@44483.4]
  assign _GEN_2145 = initBits_7 ? addrQ_7 : _GEN_2142; // @[LoadQueue.scala 308:34:@44483.4]
  assign _T_97685 = inputPriorityPorts_0_8 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44500.6]
  assign _GEN_2146 = _T_97685 ? io_addrFromLoadPorts_0 : addrQ_8; // @[LoadQueue.scala 314:36:@44504.6]
  assign _GEN_2147 = _T_97685 ? 1'h1 : addrKnown_8; // @[LoadQueue.scala 314:36:@44504.6]
  assign _GEN_2148 = initBits_8 ? 1'h0 : _GEN_2147; // @[LoadQueue.scala 308:34:@44496.4]
  assign _GEN_2149 = initBits_8 ? addrQ_8 : _GEN_2146; // @[LoadQueue.scala 308:34:@44496.4]
  assign _T_97700 = inputPriorityPorts_0_9 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44513.6]
  assign _GEN_2150 = _T_97700 ? io_addrFromLoadPorts_0 : addrQ_9; // @[LoadQueue.scala 314:36:@44517.6]
  assign _GEN_2151 = _T_97700 ? 1'h1 : addrKnown_9; // @[LoadQueue.scala 314:36:@44517.6]
  assign _GEN_2152 = initBits_9 ? 1'h0 : _GEN_2151; // @[LoadQueue.scala 308:34:@44509.4]
  assign _GEN_2153 = initBits_9 ? addrQ_9 : _GEN_2150; // @[LoadQueue.scala 308:34:@44509.4]
  assign _T_97715 = inputPriorityPorts_0_10 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44526.6]
  assign _GEN_2154 = _T_97715 ? io_addrFromLoadPorts_0 : addrQ_10; // @[LoadQueue.scala 314:36:@44530.6]
  assign _GEN_2155 = _T_97715 ? 1'h1 : addrKnown_10; // @[LoadQueue.scala 314:36:@44530.6]
  assign _GEN_2156 = initBits_10 ? 1'h0 : _GEN_2155; // @[LoadQueue.scala 308:34:@44522.4]
  assign _GEN_2157 = initBits_10 ? addrQ_10 : _GEN_2154; // @[LoadQueue.scala 308:34:@44522.4]
  assign _T_97730 = inputPriorityPorts_0_11 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44539.6]
  assign _GEN_2158 = _T_97730 ? io_addrFromLoadPorts_0 : addrQ_11; // @[LoadQueue.scala 314:36:@44543.6]
  assign _GEN_2159 = _T_97730 ? 1'h1 : addrKnown_11; // @[LoadQueue.scala 314:36:@44543.6]
  assign _GEN_2160 = initBits_11 ? 1'h0 : _GEN_2159; // @[LoadQueue.scala 308:34:@44535.4]
  assign _GEN_2161 = initBits_11 ? addrQ_11 : _GEN_2158; // @[LoadQueue.scala 308:34:@44535.4]
  assign _T_97745 = inputPriorityPorts_0_12 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44552.6]
  assign _GEN_2162 = _T_97745 ? io_addrFromLoadPorts_0 : addrQ_12; // @[LoadQueue.scala 314:36:@44556.6]
  assign _GEN_2163 = _T_97745 ? 1'h1 : addrKnown_12; // @[LoadQueue.scala 314:36:@44556.6]
  assign _GEN_2164 = initBits_12 ? 1'h0 : _GEN_2163; // @[LoadQueue.scala 308:34:@44548.4]
  assign _GEN_2165 = initBits_12 ? addrQ_12 : _GEN_2162; // @[LoadQueue.scala 308:34:@44548.4]
  assign _T_97760 = inputPriorityPorts_0_13 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44565.6]
  assign _GEN_2166 = _T_97760 ? io_addrFromLoadPorts_0 : addrQ_13; // @[LoadQueue.scala 314:36:@44569.6]
  assign _GEN_2167 = _T_97760 ? 1'h1 : addrKnown_13; // @[LoadQueue.scala 314:36:@44569.6]
  assign _GEN_2168 = initBits_13 ? 1'h0 : _GEN_2167; // @[LoadQueue.scala 308:34:@44561.4]
  assign _GEN_2169 = initBits_13 ? addrQ_13 : _GEN_2166; // @[LoadQueue.scala 308:34:@44561.4]
  assign _T_97775 = inputPriorityPorts_0_14 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44578.6]
  assign _GEN_2170 = _T_97775 ? io_addrFromLoadPorts_0 : addrQ_14; // @[LoadQueue.scala 314:36:@44582.6]
  assign _GEN_2171 = _T_97775 ? 1'h1 : addrKnown_14; // @[LoadQueue.scala 314:36:@44582.6]
  assign _GEN_2172 = initBits_14 ? 1'h0 : _GEN_2171; // @[LoadQueue.scala 308:34:@44574.4]
  assign _GEN_2173 = initBits_14 ? addrQ_14 : _GEN_2170; // @[LoadQueue.scala 308:34:@44574.4]
  assign _T_97790 = inputPriorityPorts_0_15 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@44591.6]
  assign _GEN_2174 = _T_97790 ? io_addrFromLoadPorts_0 : addrQ_15; // @[LoadQueue.scala 314:36:@44595.6]
  assign _GEN_2175 = _T_97790 ? 1'h1 : addrKnown_15; // @[LoadQueue.scala 314:36:@44595.6]
  assign _GEN_2176 = initBits_15 ? 1'h0 : _GEN_2175; // @[LoadQueue.scala 308:34:@44587.4]
  assign _GEN_2177 = initBits_15 ? addrQ_15 : _GEN_2174; // @[LoadQueue.scala 308:34:@44587.4]
  assign _T_97825 = outputPriorityPorts_0_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@44601.4]
  assign _T_97827 = loadCompleted_0 == 1'h0; // @[LoadQueue.scala 327:34:@44602.4]
  assign _T_97828 = _T_97825 & _T_97827; // @[LoadQueue.scala 327:31:@44603.4]
  assign loadCompleting_0 = _T_97828 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44604.4]
  assign _T_97839 = outputPriorityPorts_0_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@44609.4]
  assign _T_97841 = loadCompleted_1 == 1'h0; // @[LoadQueue.scala 327:34:@44610.4]
  assign _T_97842 = _T_97839 & _T_97841; // @[LoadQueue.scala 327:31:@44611.4]
  assign loadCompleting_1 = _T_97842 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44612.4]
  assign _T_97853 = outputPriorityPorts_0_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@44617.4]
  assign _T_97855 = loadCompleted_2 == 1'h0; // @[LoadQueue.scala 327:34:@44618.4]
  assign _T_97856 = _T_97853 & _T_97855; // @[LoadQueue.scala 327:31:@44619.4]
  assign loadCompleting_2 = _T_97856 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44620.4]
  assign _T_97867 = outputPriorityPorts_0_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@44625.4]
  assign _T_97869 = loadCompleted_3 == 1'h0; // @[LoadQueue.scala 327:34:@44626.4]
  assign _T_97870 = _T_97867 & _T_97869; // @[LoadQueue.scala 327:31:@44627.4]
  assign loadCompleting_3 = _T_97870 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44628.4]
  assign _T_97881 = outputPriorityPorts_0_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@44633.4]
  assign _T_97883 = loadCompleted_4 == 1'h0; // @[LoadQueue.scala 327:34:@44634.4]
  assign _T_97884 = _T_97881 & _T_97883; // @[LoadQueue.scala 327:31:@44635.4]
  assign loadCompleting_4 = _T_97884 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44636.4]
  assign _T_97895 = outputPriorityPorts_0_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@44641.4]
  assign _T_97897 = loadCompleted_5 == 1'h0; // @[LoadQueue.scala 327:34:@44642.4]
  assign _T_97898 = _T_97895 & _T_97897; // @[LoadQueue.scala 327:31:@44643.4]
  assign loadCompleting_5 = _T_97898 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44644.4]
  assign _T_97909 = outputPriorityPorts_0_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@44649.4]
  assign _T_97911 = loadCompleted_6 == 1'h0; // @[LoadQueue.scala 327:34:@44650.4]
  assign _T_97912 = _T_97909 & _T_97911; // @[LoadQueue.scala 327:31:@44651.4]
  assign loadCompleting_6 = _T_97912 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44652.4]
  assign _T_97923 = outputPriorityPorts_0_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@44657.4]
  assign _T_97925 = loadCompleted_7 == 1'h0; // @[LoadQueue.scala 327:34:@44658.4]
  assign _T_97926 = _T_97923 & _T_97925; // @[LoadQueue.scala 327:31:@44659.4]
  assign loadCompleting_7 = _T_97926 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44660.4]
  assign _T_97937 = outputPriorityPorts_0_8 & dataKnown_8; // @[LoadQueue.scala 326:108:@44665.4]
  assign _T_97939 = loadCompleted_8 == 1'h0; // @[LoadQueue.scala 327:34:@44666.4]
  assign _T_97940 = _T_97937 & _T_97939; // @[LoadQueue.scala 327:31:@44667.4]
  assign loadCompleting_8 = _T_97940 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44668.4]
  assign _T_97951 = outputPriorityPorts_0_9 & dataKnown_9; // @[LoadQueue.scala 326:108:@44673.4]
  assign _T_97953 = loadCompleted_9 == 1'h0; // @[LoadQueue.scala 327:34:@44674.4]
  assign _T_97954 = _T_97951 & _T_97953; // @[LoadQueue.scala 327:31:@44675.4]
  assign loadCompleting_9 = _T_97954 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44676.4]
  assign _T_97965 = outputPriorityPorts_0_10 & dataKnown_10; // @[LoadQueue.scala 326:108:@44681.4]
  assign _T_97967 = loadCompleted_10 == 1'h0; // @[LoadQueue.scala 327:34:@44682.4]
  assign _T_97968 = _T_97965 & _T_97967; // @[LoadQueue.scala 327:31:@44683.4]
  assign loadCompleting_10 = _T_97968 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44684.4]
  assign _T_97979 = outputPriorityPorts_0_11 & dataKnown_11; // @[LoadQueue.scala 326:108:@44689.4]
  assign _T_97981 = loadCompleted_11 == 1'h0; // @[LoadQueue.scala 327:34:@44690.4]
  assign _T_97982 = _T_97979 & _T_97981; // @[LoadQueue.scala 327:31:@44691.4]
  assign loadCompleting_11 = _T_97982 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44692.4]
  assign _T_97993 = outputPriorityPorts_0_12 & dataKnown_12; // @[LoadQueue.scala 326:108:@44697.4]
  assign _T_97995 = loadCompleted_12 == 1'h0; // @[LoadQueue.scala 327:34:@44698.4]
  assign _T_97996 = _T_97993 & _T_97995; // @[LoadQueue.scala 327:31:@44699.4]
  assign loadCompleting_12 = _T_97996 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44700.4]
  assign _T_98007 = outputPriorityPorts_0_13 & dataKnown_13; // @[LoadQueue.scala 326:108:@44705.4]
  assign _T_98009 = loadCompleted_13 == 1'h0; // @[LoadQueue.scala 327:34:@44706.4]
  assign _T_98010 = _T_98007 & _T_98009; // @[LoadQueue.scala 327:31:@44707.4]
  assign loadCompleting_13 = _T_98010 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44708.4]
  assign _T_98021 = outputPriorityPorts_0_14 & dataKnown_14; // @[LoadQueue.scala 326:108:@44713.4]
  assign _T_98023 = loadCompleted_14 == 1'h0; // @[LoadQueue.scala 327:34:@44714.4]
  assign _T_98024 = _T_98021 & _T_98023; // @[LoadQueue.scala 327:31:@44715.4]
  assign loadCompleting_14 = _T_98024 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44716.4]
  assign _T_98035 = outputPriorityPorts_0_15 & dataKnown_15; // @[LoadQueue.scala 326:108:@44721.4]
  assign _T_98037 = loadCompleted_15 == 1'h0; // @[LoadQueue.scala 327:34:@44722.4]
  assign _T_98038 = _T_98035 & _T_98037; // @[LoadQueue.scala 327:31:@44723.4]
  assign loadCompleting_15 = _T_98038 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@44724.4]
  assign _GEN_2178 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[LoadQueue.scala 337:46:@44733.6]
  assign _GEN_2179 = initBits_0 ? 1'h0 : _GEN_2178; // @[LoadQueue.scala 335:34:@44729.4]
  assign _GEN_2180 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[LoadQueue.scala 337:46:@44740.6]
  assign _GEN_2181 = initBits_1 ? 1'h0 : _GEN_2180; // @[LoadQueue.scala 335:34:@44736.4]
  assign _GEN_2182 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[LoadQueue.scala 337:46:@44747.6]
  assign _GEN_2183 = initBits_2 ? 1'h0 : _GEN_2182; // @[LoadQueue.scala 335:34:@44743.4]
  assign _GEN_2184 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[LoadQueue.scala 337:46:@44754.6]
  assign _GEN_2185 = initBits_3 ? 1'h0 : _GEN_2184; // @[LoadQueue.scala 335:34:@44750.4]
  assign _GEN_2186 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[LoadQueue.scala 337:46:@44761.6]
  assign _GEN_2187 = initBits_4 ? 1'h0 : _GEN_2186; // @[LoadQueue.scala 335:34:@44757.4]
  assign _GEN_2188 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[LoadQueue.scala 337:46:@44768.6]
  assign _GEN_2189 = initBits_5 ? 1'h0 : _GEN_2188; // @[LoadQueue.scala 335:34:@44764.4]
  assign _GEN_2190 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[LoadQueue.scala 337:46:@44775.6]
  assign _GEN_2191 = initBits_6 ? 1'h0 : _GEN_2190; // @[LoadQueue.scala 335:34:@44771.4]
  assign _GEN_2192 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[LoadQueue.scala 337:46:@44782.6]
  assign _GEN_2193 = initBits_7 ? 1'h0 : _GEN_2192; // @[LoadQueue.scala 335:34:@44778.4]
  assign _GEN_2194 = loadCompleting_8 ? 1'h1 : loadCompleted_8; // @[LoadQueue.scala 337:46:@44789.6]
  assign _GEN_2195 = initBits_8 ? 1'h0 : _GEN_2194; // @[LoadQueue.scala 335:34:@44785.4]
  assign _GEN_2196 = loadCompleting_9 ? 1'h1 : loadCompleted_9; // @[LoadQueue.scala 337:46:@44796.6]
  assign _GEN_2197 = initBits_9 ? 1'h0 : _GEN_2196; // @[LoadQueue.scala 335:34:@44792.4]
  assign _GEN_2198 = loadCompleting_10 ? 1'h1 : loadCompleted_10; // @[LoadQueue.scala 337:46:@44803.6]
  assign _GEN_2199 = initBits_10 ? 1'h0 : _GEN_2198; // @[LoadQueue.scala 335:34:@44799.4]
  assign _GEN_2200 = loadCompleting_11 ? 1'h1 : loadCompleted_11; // @[LoadQueue.scala 337:46:@44810.6]
  assign _GEN_2201 = initBits_11 ? 1'h0 : _GEN_2200; // @[LoadQueue.scala 335:34:@44806.4]
  assign _GEN_2202 = loadCompleting_12 ? 1'h1 : loadCompleted_12; // @[LoadQueue.scala 337:46:@44817.6]
  assign _GEN_2203 = initBits_12 ? 1'h0 : _GEN_2202; // @[LoadQueue.scala 335:34:@44813.4]
  assign _GEN_2204 = loadCompleting_13 ? 1'h1 : loadCompleted_13; // @[LoadQueue.scala 337:46:@44824.6]
  assign _GEN_2205 = initBits_13 ? 1'h0 : _GEN_2204; // @[LoadQueue.scala 335:34:@44820.4]
  assign _GEN_2206 = loadCompleting_14 ? 1'h1 : loadCompleted_14; // @[LoadQueue.scala 337:46:@44831.6]
  assign _GEN_2207 = initBits_14 ? 1'h0 : _GEN_2206; // @[LoadQueue.scala 335:34:@44827.4]
  assign _GEN_2208 = loadCompleting_15 ? 1'h1 : loadCompleted_15; // @[LoadQueue.scala 337:46:@44838.6]
  assign _GEN_2209 = initBits_15 ? 1'h0 : _GEN_2208; // @[LoadQueue.scala 335:34:@44834.4]
  assign _T_98169 = _T_97828 | _T_97842; // @[LoadQueue.scala 348:24:@44907.4]
  assign _T_98170 = _T_98169 | _T_97856; // @[LoadQueue.scala 348:24:@44908.4]
  assign _T_98171 = _T_98170 | _T_97870; // @[LoadQueue.scala 348:24:@44909.4]
  assign _T_98172 = _T_98171 | _T_97884; // @[LoadQueue.scala 348:24:@44910.4]
  assign _T_98173 = _T_98172 | _T_97898; // @[LoadQueue.scala 348:24:@44911.4]
  assign _T_98174 = _T_98173 | _T_97912; // @[LoadQueue.scala 348:24:@44912.4]
  assign _T_98175 = _T_98174 | _T_97926; // @[LoadQueue.scala 348:24:@44913.4]
  assign _T_98176 = _T_98175 | _T_97940; // @[LoadQueue.scala 348:24:@44914.4]
  assign _T_98177 = _T_98176 | _T_97954; // @[LoadQueue.scala 348:24:@44915.4]
  assign _T_98178 = _T_98177 | _T_97968; // @[LoadQueue.scala 348:24:@44916.4]
  assign _T_98179 = _T_98178 | _T_97982; // @[LoadQueue.scala 348:24:@44917.4]
  assign _T_98180 = _T_98179 | _T_97996; // @[LoadQueue.scala 348:24:@44918.4]
  assign _T_98181 = _T_98180 | _T_98010; // @[LoadQueue.scala 348:24:@44919.4]
  assign _T_98182 = _T_98181 | _T_98024; // @[LoadQueue.scala 348:24:@44920.4]
  assign _T_98183 = _T_98182 | _T_98038; // @[LoadQueue.scala 348:24:@44921.4]
  assign _T_98200 = _T_98024 ? 4'he : 4'hf; // @[Mux.scala 31:69:@44923.6]
  assign _T_98201 = _T_98010 ? 4'hd : _T_98200; // @[Mux.scala 31:69:@44924.6]
  assign _T_98202 = _T_97996 ? 4'hc : _T_98201; // @[Mux.scala 31:69:@44925.6]
  assign _T_98203 = _T_97982 ? 4'hb : _T_98202; // @[Mux.scala 31:69:@44926.6]
  assign _T_98204 = _T_97968 ? 4'ha : _T_98203; // @[Mux.scala 31:69:@44927.6]
  assign _T_98205 = _T_97954 ? 4'h9 : _T_98204; // @[Mux.scala 31:69:@44928.6]
  assign _T_98206 = _T_97940 ? 4'h8 : _T_98205; // @[Mux.scala 31:69:@44929.6]
  assign _T_98207 = _T_97926 ? 4'h7 : _T_98206; // @[Mux.scala 31:69:@44930.6]
  assign _T_98208 = _T_97912 ? 4'h6 : _T_98207; // @[Mux.scala 31:69:@44931.6]
  assign _T_98209 = _T_97898 ? 4'h5 : _T_98208; // @[Mux.scala 31:69:@44932.6]
  assign _T_98210 = _T_97884 ? 4'h4 : _T_98209; // @[Mux.scala 31:69:@44933.6]
  assign _T_98211 = _T_97870 ? 4'h3 : _T_98210; // @[Mux.scala 31:69:@44934.6]
  assign _T_98212 = _T_97856 ? 4'h2 : _T_98211; // @[Mux.scala 31:69:@44935.6]
  assign _T_98213 = _T_97842 ? 4'h1 : _T_98212; // @[Mux.scala 31:69:@44936.6]
  assign _T_98214 = _T_97828 ? 4'h0 : _T_98213; // @[Mux.scala 31:69:@44937.6]
  assign _GEN_2211 = 4'h1 == _T_98214 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2212 = 4'h2 == _T_98214 ? dataQ_2 : _GEN_2211; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2213 = 4'h3 == _T_98214 ? dataQ_3 : _GEN_2212; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2214 = 4'h4 == _T_98214 ? dataQ_4 : _GEN_2213; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2215 = 4'h5 == _T_98214 ? dataQ_5 : _GEN_2214; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2216 = 4'h6 == _T_98214 ? dataQ_6 : _GEN_2215; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2217 = 4'h7 == _T_98214 ? dataQ_7 : _GEN_2216; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2218 = 4'h8 == _T_98214 ? dataQ_8 : _GEN_2217; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2219 = 4'h9 == _T_98214 ? dataQ_9 : _GEN_2218; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2220 = 4'ha == _T_98214 ? dataQ_10 : _GEN_2219; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2221 = 4'hb == _T_98214 ? dataQ_11 : _GEN_2220; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2222 = 4'hc == _T_98214 ? dataQ_12 : _GEN_2221; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2223 = 4'hd == _T_98214 ? dataQ_13 : _GEN_2222; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2224 = 4'he == _T_98214 ? dataQ_14 : _GEN_2223; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2225 = 4'hf == _T_98214 ? dataQ_15 : _GEN_2224; // @[LoadQueue.scala 349:37:@44938.6]
  assign _GEN_2229 = 4'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2230 = 4'h2 == head ? loadCompleted_2 : _GEN_2229; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2231 = 4'h3 == head ? loadCompleted_3 : _GEN_2230; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2232 = 4'h4 == head ? loadCompleted_4 : _GEN_2231; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2233 = 4'h5 == head ? loadCompleted_5 : _GEN_2232; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2234 = 4'h6 == head ? loadCompleted_6 : _GEN_2233; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2235 = 4'h7 == head ? loadCompleted_7 : _GEN_2234; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2236 = 4'h8 == head ? loadCompleted_8 : _GEN_2235; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2237 = 4'h9 == head ? loadCompleted_9 : _GEN_2236; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2238 = 4'ha == head ? loadCompleted_10 : _GEN_2237; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2239 = 4'hb == head ? loadCompleted_11 : _GEN_2238; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2240 = 4'hc == head ? loadCompleted_12 : _GEN_2239; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2241 = 4'hd == head ? loadCompleted_13 : _GEN_2240; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2242 = 4'he == head ? loadCompleted_14 : _GEN_2241; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2243 = 4'hf == head ? loadCompleted_15 : _GEN_2242; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2245 = 4'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2246 = 4'h2 == head ? loadCompleting_2 : _GEN_2245; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2247 = 4'h3 == head ? loadCompleting_3 : _GEN_2246; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2248 = 4'h4 == head ? loadCompleting_4 : _GEN_2247; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2249 = 4'h5 == head ? loadCompleting_5 : _GEN_2248; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2250 = 4'h6 == head ? loadCompleting_6 : _GEN_2249; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2251 = 4'h7 == head ? loadCompleting_7 : _GEN_2250; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2252 = 4'h8 == head ? loadCompleting_8 : _GEN_2251; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2253 = 4'h9 == head ? loadCompleting_9 : _GEN_2252; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2254 = 4'ha == head ? loadCompleting_10 : _GEN_2253; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2255 = 4'hb == head ? loadCompleting_11 : _GEN_2254; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2256 = 4'hc == head ? loadCompleting_12 : _GEN_2255; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2257 = 4'hd == head ? loadCompleting_13 : _GEN_2256; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2258 = 4'he == head ? loadCompleting_14 : _GEN_2257; // @[LoadQueue.scala 363:29:@44945.4]
  assign _GEN_2259 = 4'hf == head ? loadCompleting_15 : _GEN_2258; // @[LoadQueue.scala 363:29:@44945.4]
  assign _T_98225 = _GEN_2243 | _GEN_2259; // @[LoadQueue.scala 363:29:@44945.4]
  assign _T_98226 = head != tail; // @[LoadQueue.scala 363:63:@44946.4]
  assign _T_98228 = io_loadEmpty == 1'h0; // @[LoadQueue.scala 363:75:@44947.4]
  assign _T_98229 = _T_98226 | _T_98228; // @[LoadQueue.scala 363:72:@44948.4]
  assign _T_98230 = _T_98225 & _T_98229; // @[LoadQueue.scala 363:54:@44949.4]
  assign _T_98233 = head + 4'h1; // @[util.scala 10:8:@44951.6]
  assign _GEN_64 = _T_98233 % 5'h10; // @[util.scala 10:14:@44952.6]
  assign _T_98234 = _GEN_64[4:0]; // @[util.scala 10:14:@44952.6]
  assign _GEN_2260 = _T_98230 ? _T_98234 : {{1'd0}, head}; // @[LoadQueue.scala 363:91:@44950.4]
  assign _GEN_2358 = {{3'd0}, io_bbNumLoads}; // @[util.scala 10:8:@44956.6]
  assign _T_98236 = tail + _GEN_2358; // @[util.scala 10:8:@44956.6]
  assign _GEN_65 = _T_98236 % 5'h10; // @[util.scala 10:14:@44957.6]
  assign _T_98237 = _GEN_65[4:0]; // @[util.scala 10:14:@44957.6]
  assign _GEN_2261 = io_bbStart ? _T_98237 : {{1'd0}, tail}; // @[LoadQueue.scala 367:20:@44955.4]
  assign _T_98239 = allocatedEntries_0 == 1'h0; // @[LoadQueue.scala 371:82:@44960.4]
  assign _T_98240 = loadCompleted_0 | _T_98239; // @[LoadQueue.scala 371:79:@44961.4]
  assign _T_98242 = allocatedEntries_1 == 1'h0; // @[LoadQueue.scala 371:82:@44962.4]
  assign _T_98243 = loadCompleted_1 | _T_98242; // @[LoadQueue.scala 371:79:@44963.4]
  assign _T_98245 = allocatedEntries_2 == 1'h0; // @[LoadQueue.scala 371:82:@44964.4]
  assign _T_98246 = loadCompleted_2 | _T_98245; // @[LoadQueue.scala 371:79:@44965.4]
  assign _T_98248 = allocatedEntries_3 == 1'h0; // @[LoadQueue.scala 371:82:@44966.4]
  assign _T_98249 = loadCompleted_3 | _T_98248; // @[LoadQueue.scala 371:79:@44967.4]
  assign _T_98251 = allocatedEntries_4 == 1'h0; // @[LoadQueue.scala 371:82:@44968.4]
  assign _T_98252 = loadCompleted_4 | _T_98251; // @[LoadQueue.scala 371:79:@44969.4]
  assign _T_98254 = allocatedEntries_5 == 1'h0; // @[LoadQueue.scala 371:82:@44970.4]
  assign _T_98255 = loadCompleted_5 | _T_98254; // @[LoadQueue.scala 371:79:@44971.4]
  assign _T_98257 = allocatedEntries_6 == 1'h0; // @[LoadQueue.scala 371:82:@44972.4]
  assign _T_98258 = loadCompleted_6 | _T_98257; // @[LoadQueue.scala 371:79:@44973.4]
  assign _T_98260 = allocatedEntries_7 == 1'h0; // @[LoadQueue.scala 371:82:@44974.4]
  assign _T_98261 = loadCompleted_7 | _T_98260; // @[LoadQueue.scala 371:79:@44975.4]
  assign _T_98263 = allocatedEntries_8 == 1'h0; // @[LoadQueue.scala 371:82:@44976.4]
  assign _T_98264 = loadCompleted_8 | _T_98263; // @[LoadQueue.scala 371:79:@44977.4]
  assign _T_98266 = allocatedEntries_9 == 1'h0; // @[LoadQueue.scala 371:82:@44978.4]
  assign _T_98267 = loadCompleted_9 | _T_98266; // @[LoadQueue.scala 371:79:@44979.4]
  assign _T_98269 = allocatedEntries_10 == 1'h0; // @[LoadQueue.scala 371:82:@44980.4]
  assign _T_98270 = loadCompleted_10 | _T_98269; // @[LoadQueue.scala 371:79:@44981.4]
  assign _T_98272 = allocatedEntries_11 == 1'h0; // @[LoadQueue.scala 371:82:@44982.4]
  assign _T_98273 = loadCompleted_11 | _T_98272; // @[LoadQueue.scala 371:79:@44983.4]
  assign _T_98275 = allocatedEntries_12 == 1'h0; // @[LoadQueue.scala 371:82:@44984.4]
  assign _T_98276 = loadCompleted_12 | _T_98275; // @[LoadQueue.scala 371:79:@44985.4]
  assign _T_98278 = allocatedEntries_13 == 1'h0; // @[LoadQueue.scala 371:82:@44986.4]
  assign _T_98279 = loadCompleted_13 | _T_98278; // @[LoadQueue.scala 371:79:@44987.4]
  assign _T_98281 = allocatedEntries_14 == 1'h0; // @[LoadQueue.scala 371:82:@44988.4]
  assign _T_98282 = loadCompleted_14 | _T_98281; // @[LoadQueue.scala 371:79:@44989.4]
  assign _T_98284 = allocatedEntries_15 == 1'h0; // @[LoadQueue.scala 371:82:@44990.4]
  assign _T_98285 = loadCompleted_15 | _T_98284; // @[LoadQueue.scala 371:79:@44991.4]
  assign _T_98310 = _T_98240 & _T_98243; // @[LoadQueue.scala 371:96:@45010.4]
  assign _T_98311 = _T_98310 & _T_98246; // @[LoadQueue.scala 371:96:@45011.4]
  assign _T_98312 = _T_98311 & _T_98249; // @[LoadQueue.scala 371:96:@45012.4]
  assign _T_98313 = _T_98312 & _T_98252; // @[LoadQueue.scala 371:96:@45013.4]
  assign _T_98314 = _T_98313 & _T_98255; // @[LoadQueue.scala 371:96:@45014.4]
  assign _T_98315 = _T_98314 & _T_98258; // @[LoadQueue.scala 371:96:@45015.4]
  assign _T_98316 = _T_98315 & _T_98261; // @[LoadQueue.scala 371:96:@45016.4]
  assign _T_98317 = _T_98316 & _T_98264; // @[LoadQueue.scala 371:96:@45017.4]
  assign _T_98318 = _T_98317 & _T_98267; // @[LoadQueue.scala 371:96:@45018.4]
  assign _T_98319 = _T_98318 & _T_98270; // @[LoadQueue.scala 371:96:@45019.4]
  assign _T_98320 = _T_98319 & _T_98273; // @[LoadQueue.scala 371:96:@45020.4]
  assign _T_98321 = _T_98320 & _T_98276; // @[LoadQueue.scala 371:96:@45021.4]
  assign _T_98322 = _T_98321 & _T_98279; // @[LoadQueue.scala 371:96:@45022.4]
  assign _T_98323 = _T_98322 & _T_98282; // @[LoadQueue.scala 371:96:@45023.4]
  assign io_loadTail = tail; // @[LoadQueue.scala 380:15:@45027.4]
  assign io_loadHead = head; // @[LoadQueue.scala 379:15:@45026.4]
  assign io_loadEmpty = _T_98323 & _T_98285; // @[LoadQueue.scala 371:16:@45025.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[LoadQueue.scala 382:19:@45044.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[LoadQueue.scala 382:19:@45045.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[LoadQueue.scala 382:19:@45046.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[LoadQueue.scala 382:19:@45047.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[LoadQueue.scala 382:19:@45048.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[LoadQueue.scala 382:19:@45049.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[LoadQueue.scala 382:19:@45050.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[LoadQueue.scala 382:19:@45051.4]
  assign io_loadAddrDone_8 = addrKnown_8; // @[LoadQueue.scala 382:19:@45052.4]
  assign io_loadAddrDone_9 = addrKnown_9; // @[LoadQueue.scala 382:19:@45053.4]
  assign io_loadAddrDone_10 = addrKnown_10; // @[LoadQueue.scala 382:19:@45054.4]
  assign io_loadAddrDone_11 = addrKnown_11; // @[LoadQueue.scala 382:19:@45055.4]
  assign io_loadAddrDone_12 = addrKnown_12; // @[LoadQueue.scala 382:19:@45056.4]
  assign io_loadAddrDone_13 = addrKnown_13; // @[LoadQueue.scala 382:19:@45057.4]
  assign io_loadAddrDone_14 = addrKnown_14; // @[LoadQueue.scala 382:19:@45058.4]
  assign io_loadAddrDone_15 = addrKnown_15; // @[LoadQueue.scala 382:19:@45059.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[LoadQueue.scala 383:19:@45060.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[LoadQueue.scala 383:19:@45061.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[LoadQueue.scala 383:19:@45062.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[LoadQueue.scala 383:19:@45063.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[LoadQueue.scala 383:19:@45064.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[LoadQueue.scala 383:19:@45065.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[LoadQueue.scala 383:19:@45066.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[LoadQueue.scala 383:19:@45067.4]
  assign io_loadDataDone_8 = dataKnown_8; // @[LoadQueue.scala 383:19:@45068.4]
  assign io_loadDataDone_9 = dataKnown_9; // @[LoadQueue.scala 383:19:@45069.4]
  assign io_loadDataDone_10 = dataKnown_10; // @[LoadQueue.scala 383:19:@45070.4]
  assign io_loadDataDone_11 = dataKnown_11; // @[LoadQueue.scala 383:19:@45071.4]
  assign io_loadDataDone_12 = dataKnown_12; // @[LoadQueue.scala 383:19:@45072.4]
  assign io_loadDataDone_13 = dataKnown_13; // @[LoadQueue.scala 383:19:@45073.4]
  assign io_loadDataDone_14 = dataKnown_14; // @[LoadQueue.scala 383:19:@45074.4]
  assign io_loadDataDone_15 = dataKnown_15; // @[LoadQueue.scala 383:19:@45075.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[LoadQueue.scala 381:20:@45028.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[LoadQueue.scala 381:20:@45029.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[LoadQueue.scala 381:20:@45030.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[LoadQueue.scala 381:20:@45031.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[LoadQueue.scala 381:20:@45032.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[LoadQueue.scala 381:20:@45033.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[LoadQueue.scala 381:20:@45034.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[LoadQueue.scala 381:20:@45035.4]
  assign io_loadAddrQueue_8 = addrQ_8; // @[LoadQueue.scala 381:20:@45036.4]
  assign io_loadAddrQueue_9 = addrQ_9; // @[LoadQueue.scala 381:20:@45037.4]
  assign io_loadAddrQueue_10 = addrQ_10; // @[LoadQueue.scala 381:20:@45038.4]
  assign io_loadAddrQueue_11 = addrQ_11; // @[LoadQueue.scala 381:20:@45039.4]
  assign io_loadAddrQueue_12 = addrQ_12; // @[LoadQueue.scala 381:20:@45040.4]
  assign io_loadAddrQueue_13 = addrQ_13; // @[LoadQueue.scala 381:20:@45041.4]
  assign io_loadAddrQueue_14 = addrQ_14; // @[LoadQueue.scala 381:20:@45042.4]
  assign io_loadAddrQueue_15 = addrQ_15; // @[LoadQueue.scala 381:20:@45043.4]
  assign io_loadPorts_0_valid = _T_98182 | _T_98038; // @[LoadQueue.scala 350:38:@44939.6 LoadQueue.scala 353:38:@44943.6]
  assign io_loadPorts_0_bits = _T_98183 ? _GEN_2225 : 32'h0; // @[LoadQueue.scala 349:37:@44938.6 LoadQueue.scala 352:37:@44942.6]
  assign io_loadAddrToMem = _T_93610 ? _GEN_2047 : 32'h0; // @[LoadQueue.scala 248:24:@41777.6 LoadQueue.scala 251:24:@41781.6]
  assign io_loadEnableToMem = _T_93609 | loadRequest_15; // @[LoadQueue.scala 246:22:@41744.4 LoadQueue.scala 249:26:@41778.6 LoadQueue.scala 252:26:@41782.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  loadCompleted_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  loadCompleted_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  loadCompleted_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  loadCompleted_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  loadCompleted_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  loadCompleted_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  loadCompleted_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  loadCompleted_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  bypassInitiated_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  bypassInitiated_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  bypassInitiated_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  bypassInitiated_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  bypassInitiated_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  bypassInitiated_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  bypassInitiated_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  bypassInitiated_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  checkBits_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  checkBits_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  checkBits_2 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  checkBits_3 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  checkBits_4 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  checkBits_5 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  checkBits_6 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  checkBits_7 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  checkBits_8 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  checkBits_9 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  checkBits_10 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  checkBits_11 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  checkBits_12 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  checkBits_13 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  checkBits_14 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  checkBits_15 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  previousStoreHead = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  conflictPReg_0_8 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  conflictPReg_0_9 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  conflictPReg_0_10 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  conflictPReg_0_11 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  conflictPReg_0_12 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  conflictPReg_0_13 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  conflictPReg_0_14 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  conflictPReg_0_15 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  conflictPReg_1_8 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  conflictPReg_1_9 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  conflictPReg_1_10 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  conflictPReg_1_11 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  conflictPReg_1_12 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  conflictPReg_1_13 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  conflictPReg_1_14 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  conflictPReg_1_15 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  conflictPReg_2_8 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  conflictPReg_2_9 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  conflictPReg_2_10 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  conflictPReg_2_11 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  conflictPReg_2_12 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  conflictPReg_2_13 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  conflictPReg_2_14 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  conflictPReg_2_15 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  conflictPReg_3_8 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  conflictPReg_3_9 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  conflictPReg_3_10 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  conflictPReg_3_11 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  conflictPReg_3_12 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  conflictPReg_3_13 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  conflictPReg_3_14 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  conflictPReg_3_15 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  conflictPReg_4_8 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  conflictPReg_4_9 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  conflictPReg_4_10 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  conflictPReg_4_11 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  conflictPReg_4_12 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  conflictPReg_4_13 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  conflictPReg_4_14 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  conflictPReg_4_15 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  conflictPReg_5_8 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  conflictPReg_5_9 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  conflictPReg_5_10 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  conflictPReg_5_11 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  conflictPReg_5_12 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  conflictPReg_5_13 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  conflictPReg_5_14 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  conflictPReg_5_15 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  conflictPReg_6_8 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  conflictPReg_6_9 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  conflictPReg_6_10 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  conflictPReg_6_11 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  conflictPReg_6_12 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  conflictPReg_6_13 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  conflictPReg_6_14 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  conflictPReg_6_15 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  conflictPReg_7_8 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  conflictPReg_7_9 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  conflictPReg_7_10 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  conflictPReg_7_11 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  conflictPReg_7_12 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  conflictPReg_7_13 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  conflictPReg_7_14 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  conflictPReg_7_15 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  conflictPReg_8_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  conflictPReg_8_1 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  conflictPReg_8_2 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  conflictPReg_8_3 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  conflictPReg_8_4 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  conflictPReg_8_5 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  conflictPReg_8_6 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  conflictPReg_8_7 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  conflictPReg_8_8 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  conflictPReg_8_9 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  conflictPReg_8_10 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  conflictPReg_8_11 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  conflictPReg_8_12 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  conflictPReg_8_13 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  conflictPReg_8_14 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  conflictPReg_8_15 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  conflictPReg_9_0 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  conflictPReg_9_1 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  conflictPReg_9_2 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  conflictPReg_9_3 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  conflictPReg_9_4 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  conflictPReg_9_5 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  conflictPReg_9_6 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  conflictPReg_9_7 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  conflictPReg_9_8 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  conflictPReg_9_9 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  conflictPReg_9_10 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  conflictPReg_9_11 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  conflictPReg_9_12 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  conflictPReg_9_13 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  conflictPReg_9_14 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  conflictPReg_9_15 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  conflictPReg_10_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  conflictPReg_10_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  conflictPReg_10_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  conflictPReg_10_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  conflictPReg_10_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  conflictPReg_10_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  conflictPReg_10_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  conflictPReg_10_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  conflictPReg_10_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  conflictPReg_10_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  conflictPReg_10_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  conflictPReg_10_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  conflictPReg_10_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  conflictPReg_10_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  conflictPReg_10_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  conflictPReg_10_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  conflictPReg_11_0 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  conflictPReg_11_1 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  conflictPReg_11_2 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  conflictPReg_11_3 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  conflictPReg_11_4 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  conflictPReg_11_5 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  conflictPReg_11_6 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  conflictPReg_11_7 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  conflictPReg_11_8 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  conflictPReg_11_9 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  conflictPReg_11_10 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  conflictPReg_11_11 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  conflictPReg_11_12 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  conflictPReg_11_13 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  conflictPReg_11_14 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  conflictPReg_11_15 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  conflictPReg_12_0 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  conflictPReg_12_1 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  conflictPReg_12_2 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  conflictPReg_12_3 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  conflictPReg_12_4 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  conflictPReg_12_5 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  conflictPReg_12_6 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  conflictPReg_12_7 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  conflictPReg_12_8 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  conflictPReg_12_9 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  conflictPReg_12_10 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  conflictPReg_12_11 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  conflictPReg_12_12 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  conflictPReg_12_13 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  conflictPReg_12_14 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  conflictPReg_12_15 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  conflictPReg_13_0 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  conflictPReg_13_1 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  conflictPReg_13_2 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  conflictPReg_13_3 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  conflictPReg_13_4 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  conflictPReg_13_5 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  conflictPReg_13_6 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  conflictPReg_13_7 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  conflictPReg_13_8 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  conflictPReg_13_9 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  conflictPReg_13_10 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  conflictPReg_13_11 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  conflictPReg_13_12 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  conflictPReg_13_13 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  conflictPReg_13_14 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  conflictPReg_13_15 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  conflictPReg_14_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  conflictPReg_14_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  conflictPReg_14_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  conflictPReg_14_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  conflictPReg_14_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  conflictPReg_14_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  conflictPReg_14_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  conflictPReg_14_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  conflictPReg_14_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  conflictPReg_14_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  conflictPReg_14_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  conflictPReg_14_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  conflictPReg_14_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  conflictPReg_14_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  conflictPReg_14_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  conflictPReg_14_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  conflictPReg_15_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  conflictPReg_15_1 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  conflictPReg_15_2 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  conflictPReg_15_3 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  conflictPReg_15_4 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  conflictPReg_15_5 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  conflictPReg_15_6 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  conflictPReg_15_7 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  conflictPReg_15_8 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  conflictPReg_15_9 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  conflictPReg_15_10 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  conflictPReg_15_11 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  conflictPReg_15_12 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  conflictPReg_15_13 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  conflictPReg_15_14 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  conflictPReg_15_15 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_8 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_9 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_10 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_11 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_12 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_13 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_14 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_15 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_8 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_9 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_10 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_11 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_12 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_13 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_14 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_15 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_8 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_9 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_10 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_11 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_12 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_13 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_14 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_15 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_8 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_9 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_10 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_11 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_12 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_13 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_14 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_15 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_8 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_9 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_10 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_11 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_12 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_13 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_14 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_15 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_8 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_9 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_10 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_11 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_12 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_13 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_14 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_15 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_8 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_9 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_10 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_11 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_12 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_13 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_14 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_15 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_8 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_9 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_10 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_11 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_12 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_13 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_14 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_15 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_0 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_1 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_2 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_3 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_4 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_5 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_6 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_7 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_8 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_9 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_10 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_11 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_12 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_13 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_14 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_15 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_0 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_1 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_2 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_3 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_4 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_5 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_6 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_7 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_8 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_9 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_10 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_11 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_12 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_13 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_14 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_15 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_0 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_1 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_2 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_3 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_4 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_5 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_6 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_7 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_8 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_9 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_10 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_11 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_12 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_13 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_14 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_15 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_0 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_1 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_2 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_3 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_4 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_5 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_6 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_7 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_8 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_9 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_10 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_11 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_12 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_13 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_14 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_15 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_0 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_1 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_2 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_3 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_4 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_5 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_6 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_7 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_8 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_9 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_10 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_11 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_12 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_13 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_14 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_15 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_0 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_1 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_2 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_3 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_4 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_5 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_6 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_7 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_8 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_9 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_10 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_11 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_12 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_13 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_14 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_15 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_0 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_1 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_2 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_3 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_4 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_5 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_6 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_7 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_8 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_9 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_10 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_11 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_12 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_13 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_14 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_15 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_0 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_1 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_2 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_3 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_4 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_5 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_6 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_7 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_8 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_9 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_10 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_11 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_12 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_13 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_14 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_15 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_8 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_9 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_10 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_11 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_12 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_13 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_14 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_15 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  shiftedStoreDataQPreg_8 = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  shiftedStoreDataQPreg_9 = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  shiftedStoreDataQPreg_10 = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  shiftedStoreDataQPreg_11 = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  shiftedStoreDataQPreg_12 = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  shiftedStoreDataQPreg_13 = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  shiftedStoreDataQPreg_14 = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  shiftedStoreDataQPreg_15 = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  addrKnownPReg_8 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  addrKnownPReg_9 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  addrKnownPReg_10 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  addrKnownPReg_11 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  addrKnownPReg_12 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  addrKnownPReg_13 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  addrKnownPReg_14 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  addrKnownPReg_15 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  dataKnownPReg_8 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  dataKnownPReg_9 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  dataKnownPReg_10 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  dataKnownPReg_11 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  dataKnownPReg_12 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  dataKnownPReg_13 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  dataKnownPReg_14 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  dataKnownPReg_15 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  prevPriorityRequest_15 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  prevPriorityRequest_14 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  prevPriorityRequest_13 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  prevPriorityRequest_12 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  prevPriorityRequest_11 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  prevPriorityRequest_10 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  prevPriorityRequest_9 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  prevPriorityRequest_8 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  prevPriorityRequest_7 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  prevPriorityRequest_6 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  prevPriorityRequest_5 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  prevPriorityRequest_4 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  prevPriorityRequest_3 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  prevPriorityRequest_2 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  prevPriorityRequest_1 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  prevPriorityRequest_0 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_2260[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_2261[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1924) begin
          offsetQ_0 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1924) begin
            offsetQ_0 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1924) begin
              offsetQ_0 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1924) begin
                offsetQ_0 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1924) begin
                  offsetQ_0 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1924) begin
                    offsetQ_0 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1924) begin
                      offsetQ_0 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1924) begin
                        offsetQ_0 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1924) begin
                          offsetQ_0 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1924) begin
                            offsetQ_0 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1924) begin
                              offsetQ_0 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1924) begin
                                offsetQ_0 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1924) begin
                                  offsetQ_0 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1924) begin
                                    offsetQ_0 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1924) begin
                                      offsetQ_0 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1942) begin
          offsetQ_1 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1942) begin
            offsetQ_1 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1942) begin
              offsetQ_1 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1942) begin
                offsetQ_1 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1942) begin
                  offsetQ_1 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1942) begin
                    offsetQ_1 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1942) begin
                      offsetQ_1 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1942) begin
                        offsetQ_1 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1942) begin
                          offsetQ_1 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1942) begin
                            offsetQ_1 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1942) begin
                              offsetQ_1 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1942) begin
                                offsetQ_1 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1942) begin
                                  offsetQ_1 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1942) begin
                                    offsetQ_1 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1942) begin
                                      offsetQ_1 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1960) begin
          offsetQ_2 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1960) begin
            offsetQ_2 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1960) begin
              offsetQ_2 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1960) begin
                offsetQ_2 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1960) begin
                  offsetQ_2 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1960) begin
                    offsetQ_2 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1960) begin
                      offsetQ_2 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1960) begin
                        offsetQ_2 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1960) begin
                          offsetQ_2 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1960) begin
                            offsetQ_2 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1960) begin
                              offsetQ_2 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1960) begin
                                offsetQ_2 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1960) begin
                                  offsetQ_2 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1960) begin
                                    offsetQ_2 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1960) begin
                                      offsetQ_2 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1978) begin
          offsetQ_3 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1978) begin
            offsetQ_3 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1978) begin
              offsetQ_3 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1978) begin
                offsetQ_3 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1978) begin
                  offsetQ_3 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1978) begin
                    offsetQ_3 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1978) begin
                      offsetQ_3 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1978) begin
                        offsetQ_3 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1978) begin
                          offsetQ_3 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1978) begin
                            offsetQ_3 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1978) begin
                              offsetQ_3 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1978) begin
                                offsetQ_3 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1978) begin
                                  offsetQ_3 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1978) begin
                                    offsetQ_3 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1978) begin
                                      offsetQ_3 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1996) begin
          offsetQ_4 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1996) begin
            offsetQ_4 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1996) begin
              offsetQ_4 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1996) begin
                offsetQ_4 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1996) begin
                  offsetQ_4 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1996) begin
                    offsetQ_4 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1996) begin
                      offsetQ_4 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1996) begin
                        offsetQ_4 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1996) begin
                          offsetQ_4 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1996) begin
                            offsetQ_4 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1996) begin
                              offsetQ_4 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1996) begin
                                offsetQ_4 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1996) begin
                                  offsetQ_4 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1996) begin
                                    offsetQ_4 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1996) begin
                                      offsetQ_4 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_2014) begin
          offsetQ_5 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2014) begin
            offsetQ_5 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2014) begin
              offsetQ_5 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2014) begin
                offsetQ_5 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2014) begin
                  offsetQ_5 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2014) begin
                    offsetQ_5 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2014) begin
                      offsetQ_5 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2014) begin
                        offsetQ_5 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2014) begin
                          offsetQ_5 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2014) begin
                            offsetQ_5 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2014) begin
                              offsetQ_5 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2014) begin
                                offsetQ_5 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2014) begin
                                  offsetQ_5 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2014) begin
                                    offsetQ_5 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2014) begin
                                      offsetQ_5 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_2032) begin
          offsetQ_6 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2032) begin
            offsetQ_6 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2032) begin
              offsetQ_6 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2032) begin
                offsetQ_6 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2032) begin
                  offsetQ_6 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2032) begin
                    offsetQ_6 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2032) begin
                      offsetQ_6 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2032) begin
                        offsetQ_6 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2032) begin
                          offsetQ_6 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2032) begin
                            offsetQ_6 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2032) begin
                              offsetQ_6 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2032) begin
                                offsetQ_6 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2032) begin
                                  offsetQ_6 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2032) begin
                                    offsetQ_6 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2032) begin
                                      offsetQ_6 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_2050) begin
          offsetQ_7 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2050) begin
            offsetQ_7 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2050) begin
              offsetQ_7 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2050) begin
                offsetQ_7 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2050) begin
                  offsetQ_7 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2050) begin
                    offsetQ_7 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2050) begin
                      offsetQ_7 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2050) begin
                        offsetQ_7 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2050) begin
                          offsetQ_7 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2050) begin
                            offsetQ_7 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2050) begin
                              offsetQ_7 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2050) begin
                                offsetQ_7 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2050) begin
                                  offsetQ_7 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2050) begin
                                    offsetQ_7 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2050) begin
                                      offsetQ_7 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_2068) begin
          offsetQ_8 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2068) begin
            offsetQ_8 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2068) begin
              offsetQ_8 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2068) begin
                offsetQ_8 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2068) begin
                  offsetQ_8 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2068) begin
                    offsetQ_8 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2068) begin
                      offsetQ_8 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2068) begin
                        offsetQ_8 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2068) begin
                          offsetQ_8 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2068) begin
                            offsetQ_8 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2068) begin
                              offsetQ_8 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2068) begin
                                offsetQ_8 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2068) begin
                                  offsetQ_8 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2068) begin
                                    offsetQ_8 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2068) begin
                                      offsetQ_8 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_2086) begin
          offsetQ_9 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2086) begin
            offsetQ_9 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2086) begin
              offsetQ_9 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2086) begin
                offsetQ_9 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2086) begin
                  offsetQ_9 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2086) begin
                    offsetQ_9 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2086) begin
                      offsetQ_9 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2086) begin
                        offsetQ_9 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2086) begin
                          offsetQ_9 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2086) begin
                            offsetQ_9 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2086) begin
                              offsetQ_9 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2086) begin
                                offsetQ_9 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2086) begin
                                  offsetQ_9 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2086) begin
                                    offsetQ_9 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2086) begin
                                      offsetQ_9 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_2104) begin
          offsetQ_10 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2104) begin
            offsetQ_10 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2104) begin
              offsetQ_10 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2104) begin
                offsetQ_10 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2104) begin
                  offsetQ_10 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2104) begin
                    offsetQ_10 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2104) begin
                      offsetQ_10 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2104) begin
                        offsetQ_10 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2104) begin
                          offsetQ_10 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2104) begin
                            offsetQ_10 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2104) begin
                              offsetQ_10 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2104) begin
                                offsetQ_10 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2104) begin
                                  offsetQ_10 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2104) begin
                                    offsetQ_10 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2104) begin
                                      offsetQ_10 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2122) begin
          offsetQ_11 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2122) begin
            offsetQ_11 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2122) begin
              offsetQ_11 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2122) begin
                offsetQ_11 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2122) begin
                  offsetQ_11 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2122) begin
                    offsetQ_11 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2122) begin
                      offsetQ_11 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2122) begin
                        offsetQ_11 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2122) begin
                          offsetQ_11 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2122) begin
                            offsetQ_11 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2122) begin
                              offsetQ_11 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2122) begin
                                offsetQ_11 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2122) begin
                                  offsetQ_11 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2122) begin
                                    offsetQ_11 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2122) begin
                                      offsetQ_11 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2140) begin
          offsetQ_12 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2140) begin
            offsetQ_12 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2140) begin
              offsetQ_12 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2140) begin
                offsetQ_12 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2140) begin
                  offsetQ_12 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2140) begin
                    offsetQ_12 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2140) begin
                      offsetQ_12 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2140) begin
                        offsetQ_12 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2140) begin
                          offsetQ_12 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2140) begin
                            offsetQ_12 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2140) begin
                              offsetQ_12 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2140) begin
                                offsetQ_12 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2140) begin
                                  offsetQ_12 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2140) begin
                                    offsetQ_12 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2140) begin
                                      offsetQ_12 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2158) begin
          offsetQ_13 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2158) begin
            offsetQ_13 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2158) begin
              offsetQ_13 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2158) begin
                offsetQ_13 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2158) begin
                  offsetQ_13 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2158) begin
                    offsetQ_13 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2158) begin
                      offsetQ_13 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2158) begin
                        offsetQ_13 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2158) begin
                          offsetQ_13 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2158) begin
                            offsetQ_13 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2158) begin
                              offsetQ_13 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2158) begin
                                offsetQ_13 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2158) begin
                                  offsetQ_13 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2158) begin
                                    offsetQ_13 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2158) begin
                                      offsetQ_13 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2176) begin
          offsetQ_14 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2176) begin
            offsetQ_14 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2176) begin
              offsetQ_14 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2176) begin
                offsetQ_14 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2176) begin
                  offsetQ_14 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2176) begin
                    offsetQ_14 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2176) begin
                      offsetQ_14 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2176) begin
                        offsetQ_14 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2176) begin
                          offsetQ_14 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2176) begin
                            offsetQ_14 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2176) begin
                              offsetQ_14 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2176) begin
                                offsetQ_14 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2176) begin
                                  offsetQ_14 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2176) begin
                                    offsetQ_14 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2176) begin
                                      offsetQ_14 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2194) begin
          offsetQ_15 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2194) begin
            offsetQ_15 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2194) begin
              offsetQ_15 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2194) begin
                offsetQ_15 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2194) begin
                  offsetQ_15 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2194) begin
                    offsetQ_15 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2194) begin
                      offsetQ_15 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2194) begin
                        offsetQ_15 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2194) begin
                          offsetQ_15 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2194) begin
                            offsetQ_15 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2194) begin
                              offsetQ_15 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2194) begin
                                offsetQ_15 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2194) begin
                                  offsetQ_15 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2194) begin
                                    offsetQ_15 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2194) begin
                                      offsetQ_15 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_97565) begin
          addrQ_0 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_97580) begin
          addrQ_1 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_97595) begin
          addrQ_2 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_97610) begin
          addrQ_3 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_97625) begin
          addrQ_4 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_97640) begin
          addrQ_5 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_97655) begin
          addrQ_6 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_97670) begin
          addrQ_7 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_97685) begin
          addrQ_8 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_97700) begin
          addrQ_9 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_97715) begin
          addrQ_10 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_97730) begin
          addrQ_11 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_97745) begin
          addrQ_12 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_97760) begin
          addrQ_13 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_97775) begin
          addrQ_14 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_97790) begin
          addrQ_15 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_88298) begin
          if (4'hf == _T_88281) begin
            dataQ_0 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88281) begin
              dataQ_0 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88281) begin
                dataQ_0 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88281) begin
                  dataQ_0 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88281) begin
                    dataQ_0 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88281) begin
                      dataQ_0 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88281) begin
                        dataQ_0 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88281) begin
                          dataQ_0 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88281) begin
                            dataQ_0 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88281) begin
                              dataQ_0 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88281) begin
                                dataQ_0 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88281) begin
                                  dataQ_0 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88281) begin
                                    dataQ_0 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88281) begin
                                      dataQ_0 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88281) begin
                                        dataQ_0 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_0 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_0) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_88434) begin
          if (4'hf == _T_88417) begin
            dataQ_1 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88417) begin
              dataQ_1 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88417) begin
                dataQ_1 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88417) begin
                  dataQ_1 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88417) begin
                    dataQ_1 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88417) begin
                      dataQ_1 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88417) begin
                        dataQ_1 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88417) begin
                          dataQ_1 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88417) begin
                            dataQ_1 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88417) begin
                              dataQ_1 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88417) begin
                                dataQ_1 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88417) begin
                                  dataQ_1 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88417) begin
                                    dataQ_1 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88417) begin
                                      dataQ_1 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88417) begin
                                        dataQ_1 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_1 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_1) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_88570) begin
          if (4'hf == _T_88553) begin
            dataQ_2 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88553) begin
              dataQ_2 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88553) begin
                dataQ_2 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88553) begin
                  dataQ_2 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88553) begin
                    dataQ_2 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88553) begin
                      dataQ_2 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88553) begin
                        dataQ_2 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88553) begin
                          dataQ_2 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88553) begin
                            dataQ_2 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88553) begin
                              dataQ_2 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88553) begin
                                dataQ_2 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88553) begin
                                  dataQ_2 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88553) begin
                                    dataQ_2 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88553) begin
                                      dataQ_2 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88553) begin
                                        dataQ_2 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_2 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_2) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_88706) begin
          if (4'hf == _T_88689) begin
            dataQ_3 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88689) begin
              dataQ_3 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88689) begin
                dataQ_3 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88689) begin
                  dataQ_3 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88689) begin
                    dataQ_3 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88689) begin
                      dataQ_3 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88689) begin
                        dataQ_3 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88689) begin
                          dataQ_3 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88689) begin
                            dataQ_3 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88689) begin
                              dataQ_3 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88689) begin
                                dataQ_3 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88689) begin
                                  dataQ_3 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88689) begin
                                    dataQ_3 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88689) begin
                                      dataQ_3 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88689) begin
                                        dataQ_3 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_3 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_3) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_88842) begin
          if (4'hf == _T_88825) begin
            dataQ_4 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88825) begin
              dataQ_4 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88825) begin
                dataQ_4 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88825) begin
                  dataQ_4 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88825) begin
                    dataQ_4 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88825) begin
                      dataQ_4 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88825) begin
                        dataQ_4 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88825) begin
                          dataQ_4 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88825) begin
                            dataQ_4 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88825) begin
                              dataQ_4 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88825) begin
                                dataQ_4 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88825) begin
                                  dataQ_4 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88825) begin
                                    dataQ_4 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88825) begin
                                      dataQ_4 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88825) begin
                                        dataQ_4 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_4 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_4) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_88978) begin
          if (4'hf == _T_88961) begin
            dataQ_5 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88961) begin
              dataQ_5 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88961) begin
                dataQ_5 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88961) begin
                  dataQ_5 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88961) begin
                    dataQ_5 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88961) begin
                      dataQ_5 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88961) begin
                        dataQ_5 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88961) begin
                          dataQ_5 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88961) begin
                            dataQ_5 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88961) begin
                              dataQ_5 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88961) begin
                                dataQ_5 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88961) begin
                                  dataQ_5 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88961) begin
                                    dataQ_5 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88961) begin
                                      dataQ_5 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88961) begin
                                        dataQ_5 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_5 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_5) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_89114) begin
          if (4'hf == _T_89097) begin
            dataQ_6 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89097) begin
              dataQ_6 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89097) begin
                dataQ_6 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89097) begin
                  dataQ_6 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89097) begin
                    dataQ_6 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89097) begin
                      dataQ_6 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89097) begin
                        dataQ_6 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89097) begin
                          dataQ_6 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89097) begin
                            dataQ_6 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89097) begin
                              dataQ_6 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89097) begin
                                dataQ_6 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89097) begin
                                  dataQ_6 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89097) begin
                                    dataQ_6 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89097) begin
                                      dataQ_6 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89097) begin
                                        dataQ_6 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_6 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_6) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_89250) begin
          if (4'hf == _T_89233) begin
            dataQ_7 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89233) begin
              dataQ_7 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89233) begin
                dataQ_7 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89233) begin
                  dataQ_7 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89233) begin
                    dataQ_7 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89233) begin
                      dataQ_7 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89233) begin
                        dataQ_7 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89233) begin
                          dataQ_7 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89233) begin
                            dataQ_7 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89233) begin
                              dataQ_7 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89233) begin
                                dataQ_7 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89233) begin
                                  dataQ_7 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89233) begin
                                    dataQ_7 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89233) begin
                                      dataQ_7 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89233) begin
                                        dataQ_7 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_7 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_7) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (bypassRequest_8) begin
        if (_T_89386) begin
          if (4'hf == _T_89369) begin
            dataQ_8 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89369) begin
              dataQ_8 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89369) begin
                dataQ_8 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89369) begin
                  dataQ_8 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89369) begin
                    dataQ_8 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89369) begin
                      dataQ_8 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89369) begin
                        dataQ_8 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89369) begin
                          dataQ_8 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89369) begin
                            dataQ_8 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89369) begin
                              dataQ_8 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89369) begin
                                dataQ_8 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89369) begin
                                  dataQ_8 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89369) begin
                                    dataQ_8 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89369) begin
                                      dataQ_8 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89369) begin
                                        dataQ_8 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_8 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_8 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_8) begin
          dataQ_8 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (bypassRequest_9) begin
        if (_T_89522) begin
          if (4'hf == _T_89505) begin
            dataQ_9 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89505) begin
              dataQ_9 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89505) begin
                dataQ_9 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89505) begin
                  dataQ_9 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89505) begin
                    dataQ_9 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89505) begin
                      dataQ_9 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89505) begin
                        dataQ_9 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89505) begin
                          dataQ_9 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89505) begin
                            dataQ_9 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89505) begin
                              dataQ_9 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89505) begin
                                dataQ_9 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89505) begin
                                  dataQ_9 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89505) begin
                                    dataQ_9 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89505) begin
                                      dataQ_9 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89505) begin
                                        dataQ_9 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_9 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_9 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_9) begin
          dataQ_9 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (bypassRequest_10) begin
        if (_T_89658) begin
          if (4'hf == _T_89641) begin
            dataQ_10 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89641) begin
              dataQ_10 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89641) begin
                dataQ_10 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89641) begin
                  dataQ_10 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89641) begin
                    dataQ_10 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89641) begin
                      dataQ_10 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89641) begin
                        dataQ_10 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89641) begin
                          dataQ_10 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89641) begin
                            dataQ_10 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89641) begin
                              dataQ_10 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89641) begin
                                dataQ_10 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89641) begin
                                  dataQ_10 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89641) begin
                                    dataQ_10 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89641) begin
                                      dataQ_10 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89641) begin
                                        dataQ_10 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_10 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_10 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_10) begin
          dataQ_10 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (bypassRequest_11) begin
        if (_T_89794) begin
          if (4'hf == _T_89777) begin
            dataQ_11 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89777) begin
              dataQ_11 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89777) begin
                dataQ_11 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89777) begin
                  dataQ_11 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89777) begin
                    dataQ_11 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89777) begin
                      dataQ_11 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89777) begin
                        dataQ_11 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89777) begin
                          dataQ_11 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89777) begin
                            dataQ_11 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89777) begin
                              dataQ_11 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89777) begin
                                dataQ_11 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89777) begin
                                  dataQ_11 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89777) begin
                                    dataQ_11 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89777) begin
                                      dataQ_11 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89777) begin
                                        dataQ_11 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_11 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_11 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_11) begin
          dataQ_11 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (bypassRequest_12) begin
        if (_T_89930) begin
          if (4'hf == _T_89913) begin
            dataQ_12 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89913) begin
              dataQ_12 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89913) begin
                dataQ_12 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89913) begin
                  dataQ_12 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89913) begin
                    dataQ_12 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89913) begin
                      dataQ_12 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89913) begin
                        dataQ_12 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89913) begin
                          dataQ_12 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89913) begin
                            dataQ_12 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89913) begin
                              dataQ_12 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89913) begin
                                dataQ_12 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89913) begin
                                  dataQ_12 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89913) begin
                                    dataQ_12 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89913) begin
                                      dataQ_12 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89913) begin
                                        dataQ_12 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_12 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_12 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_12) begin
          dataQ_12 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (bypassRequest_13) begin
        if (_T_90066) begin
          if (4'hf == _T_90049) begin
            dataQ_13 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90049) begin
              dataQ_13 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90049) begin
                dataQ_13 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90049) begin
                  dataQ_13 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90049) begin
                    dataQ_13 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90049) begin
                      dataQ_13 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90049) begin
                        dataQ_13 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90049) begin
                          dataQ_13 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90049) begin
                            dataQ_13 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90049) begin
                              dataQ_13 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90049) begin
                                dataQ_13 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90049) begin
                                  dataQ_13 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90049) begin
                                    dataQ_13 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90049) begin
                                      dataQ_13 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90049) begin
                                        dataQ_13 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_13 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_13 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_13) begin
          dataQ_13 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (bypassRequest_14) begin
        if (_T_90202) begin
          if (4'hf == _T_90185) begin
            dataQ_14 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90185) begin
              dataQ_14 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90185) begin
                dataQ_14 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90185) begin
                  dataQ_14 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90185) begin
                    dataQ_14 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90185) begin
                      dataQ_14 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90185) begin
                        dataQ_14 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90185) begin
                          dataQ_14 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90185) begin
                            dataQ_14 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90185) begin
                              dataQ_14 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90185) begin
                                dataQ_14 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90185) begin
                                  dataQ_14 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90185) begin
                                    dataQ_14 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90185) begin
                                      dataQ_14 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90185) begin
                                        dataQ_14 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_14 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_14 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_14) begin
          dataQ_14 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (bypassRequest_15) begin
        if (_T_90338) begin
          if (4'hf == _T_90321) begin
            dataQ_15 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90321) begin
              dataQ_15 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90321) begin
                dataQ_15 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90321) begin
                  dataQ_15 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90321) begin
                    dataQ_15 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90321) begin
                      dataQ_15 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90321) begin
                        dataQ_15 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90321) begin
                          dataQ_15 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90321) begin
                            dataQ_15 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90321) begin
                              dataQ_15 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90321) begin
                                dataQ_15 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90321) begin
                                  dataQ_15 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90321) begin
                                    dataQ_15 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90321) begin
                                      dataQ_15 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90321) begin
                                        dataQ_15 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_15 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_15 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_15) begin
          dataQ_15 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_97565) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_97580) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_97595) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_97610) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_97625) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_97640) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_97655) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_97670) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_97685) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_97700) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_97715) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_97730) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_97745) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_97760) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_97775) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_97790) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_93649) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_93652) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_93655) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_93658) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_93661) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_93664) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_93667) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_93670) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_93673) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_93676) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_93679) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_93682) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_93685) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_93688) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_93691) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_93694) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        loadCompleted_8 <= 1'h0;
      end else begin
        if (loadCompleting_8) begin
          loadCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        loadCompleted_9 <= 1'h0;
      end else begin
        if (loadCompleting_9) begin
          loadCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        loadCompleted_10 <= 1'h0;
      end else begin
        if (loadCompleting_10) begin
          loadCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        loadCompleted_11 <= 1'h0;
      end else begin
        if (loadCompleting_11) begin
          loadCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        loadCompleted_12 <= 1'h0;
      end else begin
        if (loadCompleting_12) begin
          loadCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        loadCompleted_13 <= 1'h0;
      end else begin
        if (loadCompleting_13) begin
          loadCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        loadCompleted_14 <= 1'h0;
      end else begin
        if (loadCompleting_14) begin
          loadCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        loadCompleted_15 <= 1'h0;
      end else begin
        if (loadCompleting_15) begin
          loadCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1878;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1879;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1880;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1881;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1882;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1883;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1884;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1885;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1886;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1887;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1888;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1889;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1890;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1891;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1892;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1893;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        bypassInitiated_8 <= 1'h0;
      end else begin
        if (bypassRequest_8) begin
          bypassInitiated_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        bypassInitiated_9 <= 1'h0;
      end else begin
        if (bypassRequest_9) begin
          bypassInitiated_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        bypassInitiated_10 <= 1'h0;
      end else begin
        if (bypassRequest_10) begin
          bypassInitiated_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        bypassInitiated_11 <= 1'h0;
      end else begin
        if (bypassRequest_11) begin
          bypassInitiated_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        bypassInitiated_12 <= 1'h0;
      end else begin
        if (bypassRequest_12) begin
          bypassInitiated_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        bypassInitiated_13 <= 1'h0;
      end else begin
        if (bypassRequest_13) begin
          bypassInitiated_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        bypassInitiated_14 <= 1'h0;
      end else begin
        if (bypassRequest_14) begin
          bypassInitiated_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        bypassInitiated_15 <= 1'h0;
      end else begin
        if (bypassRequest_15) begin
          bypassInitiated_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2221;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2225) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2233) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2251;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2255) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2263) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2281;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2285) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2293) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2311;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2315) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2323) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2341;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2345) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2353) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2371;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2375) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2383) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2401;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2405) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2413) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2431;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2435) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2443) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2461;
      end else begin
        if (io_storeEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2465) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2473) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2491;
      end else begin
        if (io_storeEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2495) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2503) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2521;
      end else begin
        if (io_storeEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2525) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2533) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2551;
      end else begin
        if (io_storeEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2555) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2563) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2581;
      end else begin
        if (io_storeEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2585) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2593) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2611;
      end else begin
        if (io_storeEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2615) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2623) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2641;
      end else begin
        if (io_storeEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2645) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2653) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2671;
      end else begin
        if (io_storeEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2675) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2683) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_18282[0];
    conflictPReg_0_1 <= _T_18282[1];
    conflictPReg_0_2 <= _T_18282[2];
    conflictPReg_0_3 <= _T_18282[3];
    conflictPReg_0_4 <= _T_18282[4];
    conflictPReg_0_5 <= _T_18282[5];
    conflictPReg_0_6 <= _T_18282[6];
    conflictPReg_0_7 <= _T_18282[7];
    conflictPReg_0_8 <= _T_18282[8];
    conflictPReg_0_9 <= _T_18282[9];
    conflictPReg_0_10 <= _T_18282[10];
    conflictPReg_0_11 <= _T_18282[11];
    conflictPReg_0_12 <= _T_18282[12];
    conflictPReg_0_13 <= _T_18282[13];
    conflictPReg_0_14 <= _T_18282[14];
    conflictPReg_0_15 <= _T_18282[15];
    conflictPReg_1_0 <= _T_19140[0];
    conflictPReg_1_1 <= _T_19140[1];
    conflictPReg_1_2 <= _T_19140[2];
    conflictPReg_1_3 <= _T_19140[3];
    conflictPReg_1_4 <= _T_19140[4];
    conflictPReg_1_5 <= _T_19140[5];
    conflictPReg_1_6 <= _T_19140[6];
    conflictPReg_1_7 <= _T_19140[7];
    conflictPReg_1_8 <= _T_19140[8];
    conflictPReg_1_9 <= _T_19140[9];
    conflictPReg_1_10 <= _T_19140[10];
    conflictPReg_1_11 <= _T_19140[11];
    conflictPReg_1_12 <= _T_19140[12];
    conflictPReg_1_13 <= _T_19140[13];
    conflictPReg_1_14 <= _T_19140[14];
    conflictPReg_1_15 <= _T_19140[15];
    conflictPReg_2_0 <= _T_19998[0];
    conflictPReg_2_1 <= _T_19998[1];
    conflictPReg_2_2 <= _T_19998[2];
    conflictPReg_2_3 <= _T_19998[3];
    conflictPReg_2_4 <= _T_19998[4];
    conflictPReg_2_5 <= _T_19998[5];
    conflictPReg_2_6 <= _T_19998[6];
    conflictPReg_2_7 <= _T_19998[7];
    conflictPReg_2_8 <= _T_19998[8];
    conflictPReg_2_9 <= _T_19998[9];
    conflictPReg_2_10 <= _T_19998[10];
    conflictPReg_2_11 <= _T_19998[11];
    conflictPReg_2_12 <= _T_19998[12];
    conflictPReg_2_13 <= _T_19998[13];
    conflictPReg_2_14 <= _T_19998[14];
    conflictPReg_2_15 <= _T_19998[15];
    conflictPReg_3_0 <= _T_20856[0];
    conflictPReg_3_1 <= _T_20856[1];
    conflictPReg_3_2 <= _T_20856[2];
    conflictPReg_3_3 <= _T_20856[3];
    conflictPReg_3_4 <= _T_20856[4];
    conflictPReg_3_5 <= _T_20856[5];
    conflictPReg_3_6 <= _T_20856[6];
    conflictPReg_3_7 <= _T_20856[7];
    conflictPReg_3_8 <= _T_20856[8];
    conflictPReg_3_9 <= _T_20856[9];
    conflictPReg_3_10 <= _T_20856[10];
    conflictPReg_3_11 <= _T_20856[11];
    conflictPReg_3_12 <= _T_20856[12];
    conflictPReg_3_13 <= _T_20856[13];
    conflictPReg_3_14 <= _T_20856[14];
    conflictPReg_3_15 <= _T_20856[15];
    conflictPReg_4_0 <= _T_21714[0];
    conflictPReg_4_1 <= _T_21714[1];
    conflictPReg_4_2 <= _T_21714[2];
    conflictPReg_4_3 <= _T_21714[3];
    conflictPReg_4_4 <= _T_21714[4];
    conflictPReg_4_5 <= _T_21714[5];
    conflictPReg_4_6 <= _T_21714[6];
    conflictPReg_4_7 <= _T_21714[7];
    conflictPReg_4_8 <= _T_21714[8];
    conflictPReg_4_9 <= _T_21714[9];
    conflictPReg_4_10 <= _T_21714[10];
    conflictPReg_4_11 <= _T_21714[11];
    conflictPReg_4_12 <= _T_21714[12];
    conflictPReg_4_13 <= _T_21714[13];
    conflictPReg_4_14 <= _T_21714[14];
    conflictPReg_4_15 <= _T_21714[15];
    conflictPReg_5_0 <= _T_22572[0];
    conflictPReg_5_1 <= _T_22572[1];
    conflictPReg_5_2 <= _T_22572[2];
    conflictPReg_5_3 <= _T_22572[3];
    conflictPReg_5_4 <= _T_22572[4];
    conflictPReg_5_5 <= _T_22572[5];
    conflictPReg_5_6 <= _T_22572[6];
    conflictPReg_5_7 <= _T_22572[7];
    conflictPReg_5_8 <= _T_22572[8];
    conflictPReg_5_9 <= _T_22572[9];
    conflictPReg_5_10 <= _T_22572[10];
    conflictPReg_5_11 <= _T_22572[11];
    conflictPReg_5_12 <= _T_22572[12];
    conflictPReg_5_13 <= _T_22572[13];
    conflictPReg_5_14 <= _T_22572[14];
    conflictPReg_5_15 <= _T_22572[15];
    conflictPReg_6_0 <= _T_23430[0];
    conflictPReg_6_1 <= _T_23430[1];
    conflictPReg_6_2 <= _T_23430[2];
    conflictPReg_6_3 <= _T_23430[3];
    conflictPReg_6_4 <= _T_23430[4];
    conflictPReg_6_5 <= _T_23430[5];
    conflictPReg_6_6 <= _T_23430[6];
    conflictPReg_6_7 <= _T_23430[7];
    conflictPReg_6_8 <= _T_23430[8];
    conflictPReg_6_9 <= _T_23430[9];
    conflictPReg_6_10 <= _T_23430[10];
    conflictPReg_6_11 <= _T_23430[11];
    conflictPReg_6_12 <= _T_23430[12];
    conflictPReg_6_13 <= _T_23430[13];
    conflictPReg_6_14 <= _T_23430[14];
    conflictPReg_6_15 <= _T_23430[15];
    conflictPReg_7_0 <= _T_24288[0];
    conflictPReg_7_1 <= _T_24288[1];
    conflictPReg_7_2 <= _T_24288[2];
    conflictPReg_7_3 <= _T_24288[3];
    conflictPReg_7_4 <= _T_24288[4];
    conflictPReg_7_5 <= _T_24288[5];
    conflictPReg_7_6 <= _T_24288[6];
    conflictPReg_7_7 <= _T_24288[7];
    conflictPReg_7_8 <= _T_24288[8];
    conflictPReg_7_9 <= _T_24288[9];
    conflictPReg_7_10 <= _T_24288[10];
    conflictPReg_7_11 <= _T_24288[11];
    conflictPReg_7_12 <= _T_24288[12];
    conflictPReg_7_13 <= _T_24288[13];
    conflictPReg_7_14 <= _T_24288[14];
    conflictPReg_7_15 <= _T_24288[15];
    conflictPReg_8_0 <= _T_25146[0];
    conflictPReg_8_1 <= _T_25146[1];
    conflictPReg_8_2 <= _T_25146[2];
    conflictPReg_8_3 <= _T_25146[3];
    conflictPReg_8_4 <= _T_25146[4];
    conflictPReg_8_5 <= _T_25146[5];
    conflictPReg_8_6 <= _T_25146[6];
    conflictPReg_8_7 <= _T_25146[7];
    conflictPReg_8_8 <= _T_25146[8];
    conflictPReg_8_9 <= _T_25146[9];
    conflictPReg_8_10 <= _T_25146[10];
    conflictPReg_8_11 <= _T_25146[11];
    conflictPReg_8_12 <= _T_25146[12];
    conflictPReg_8_13 <= _T_25146[13];
    conflictPReg_8_14 <= _T_25146[14];
    conflictPReg_8_15 <= _T_25146[15];
    conflictPReg_9_0 <= _T_26004[0];
    conflictPReg_9_1 <= _T_26004[1];
    conflictPReg_9_2 <= _T_26004[2];
    conflictPReg_9_3 <= _T_26004[3];
    conflictPReg_9_4 <= _T_26004[4];
    conflictPReg_9_5 <= _T_26004[5];
    conflictPReg_9_6 <= _T_26004[6];
    conflictPReg_9_7 <= _T_26004[7];
    conflictPReg_9_8 <= _T_26004[8];
    conflictPReg_9_9 <= _T_26004[9];
    conflictPReg_9_10 <= _T_26004[10];
    conflictPReg_9_11 <= _T_26004[11];
    conflictPReg_9_12 <= _T_26004[12];
    conflictPReg_9_13 <= _T_26004[13];
    conflictPReg_9_14 <= _T_26004[14];
    conflictPReg_9_15 <= _T_26004[15];
    conflictPReg_10_0 <= _T_26862[0];
    conflictPReg_10_1 <= _T_26862[1];
    conflictPReg_10_2 <= _T_26862[2];
    conflictPReg_10_3 <= _T_26862[3];
    conflictPReg_10_4 <= _T_26862[4];
    conflictPReg_10_5 <= _T_26862[5];
    conflictPReg_10_6 <= _T_26862[6];
    conflictPReg_10_7 <= _T_26862[7];
    conflictPReg_10_8 <= _T_26862[8];
    conflictPReg_10_9 <= _T_26862[9];
    conflictPReg_10_10 <= _T_26862[10];
    conflictPReg_10_11 <= _T_26862[11];
    conflictPReg_10_12 <= _T_26862[12];
    conflictPReg_10_13 <= _T_26862[13];
    conflictPReg_10_14 <= _T_26862[14];
    conflictPReg_10_15 <= _T_26862[15];
    conflictPReg_11_0 <= _T_27720[0];
    conflictPReg_11_1 <= _T_27720[1];
    conflictPReg_11_2 <= _T_27720[2];
    conflictPReg_11_3 <= _T_27720[3];
    conflictPReg_11_4 <= _T_27720[4];
    conflictPReg_11_5 <= _T_27720[5];
    conflictPReg_11_6 <= _T_27720[6];
    conflictPReg_11_7 <= _T_27720[7];
    conflictPReg_11_8 <= _T_27720[8];
    conflictPReg_11_9 <= _T_27720[9];
    conflictPReg_11_10 <= _T_27720[10];
    conflictPReg_11_11 <= _T_27720[11];
    conflictPReg_11_12 <= _T_27720[12];
    conflictPReg_11_13 <= _T_27720[13];
    conflictPReg_11_14 <= _T_27720[14];
    conflictPReg_11_15 <= _T_27720[15];
    conflictPReg_12_0 <= _T_28578[0];
    conflictPReg_12_1 <= _T_28578[1];
    conflictPReg_12_2 <= _T_28578[2];
    conflictPReg_12_3 <= _T_28578[3];
    conflictPReg_12_4 <= _T_28578[4];
    conflictPReg_12_5 <= _T_28578[5];
    conflictPReg_12_6 <= _T_28578[6];
    conflictPReg_12_7 <= _T_28578[7];
    conflictPReg_12_8 <= _T_28578[8];
    conflictPReg_12_9 <= _T_28578[9];
    conflictPReg_12_10 <= _T_28578[10];
    conflictPReg_12_11 <= _T_28578[11];
    conflictPReg_12_12 <= _T_28578[12];
    conflictPReg_12_13 <= _T_28578[13];
    conflictPReg_12_14 <= _T_28578[14];
    conflictPReg_12_15 <= _T_28578[15];
    conflictPReg_13_0 <= _T_29436[0];
    conflictPReg_13_1 <= _T_29436[1];
    conflictPReg_13_2 <= _T_29436[2];
    conflictPReg_13_3 <= _T_29436[3];
    conflictPReg_13_4 <= _T_29436[4];
    conflictPReg_13_5 <= _T_29436[5];
    conflictPReg_13_6 <= _T_29436[6];
    conflictPReg_13_7 <= _T_29436[7];
    conflictPReg_13_8 <= _T_29436[8];
    conflictPReg_13_9 <= _T_29436[9];
    conflictPReg_13_10 <= _T_29436[10];
    conflictPReg_13_11 <= _T_29436[11];
    conflictPReg_13_12 <= _T_29436[12];
    conflictPReg_13_13 <= _T_29436[13];
    conflictPReg_13_14 <= _T_29436[14];
    conflictPReg_13_15 <= _T_29436[15];
    conflictPReg_14_0 <= _T_30294[0];
    conflictPReg_14_1 <= _T_30294[1];
    conflictPReg_14_2 <= _T_30294[2];
    conflictPReg_14_3 <= _T_30294[3];
    conflictPReg_14_4 <= _T_30294[4];
    conflictPReg_14_5 <= _T_30294[5];
    conflictPReg_14_6 <= _T_30294[6];
    conflictPReg_14_7 <= _T_30294[7];
    conflictPReg_14_8 <= _T_30294[8];
    conflictPReg_14_9 <= _T_30294[9];
    conflictPReg_14_10 <= _T_30294[10];
    conflictPReg_14_11 <= _T_30294[11];
    conflictPReg_14_12 <= _T_30294[12];
    conflictPReg_14_13 <= _T_30294[13];
    conflictPReg_14_14 <= _T_30294[14];
    conflictPReg_14_15 <= _T_30294[15];
    conflictPReg_15_0 <= _T_31152[0];
    conflictPReg_15_1 <= _T_31152[1];
    conflictPReg_15_2 <= _T_31152[2];
    conflictPReg_15_3 <= _T_31152[3];
    conflictPReg_15_4 <= _T_31152[4];
    conflictPReg_15_5 <= _T_31152[5];
    conflictPReg_15_6 <= _T_31152[6];
    conflictPReg_15_7 <= _T_31152[7];
    conflictPReg_15_8 <= _T_31152[8];
    conflictPReg_15_9 <= _T_31152[9];
    conflictPReg_15_10 <= _T_31152[10];
    conflictPReg_15_11 <= _T_31152[11];
    conflictPReg_15_12 <= _T_31152[12];
    conflictPReg_15_13 <= _T_31152[13];
    conflictPReg_15_14 <= _T_31152[14];
    conflictPReg_15_15 <= _T_31152[15];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_52606[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_52606[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_52606[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_52606[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_52606[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_52606[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_52606[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_52606[7];
    storeAddrNotKnownFlagsPReg_0_8 <= _T_52606[8];
    storeAddrNotKnownFlagsPReg_0_9 <= _T_52606[9];
    storeAddrNotKnownFlagsPReg_0_10 <= _T_52606[10];
    storeAddrNotKnownFlagsPReg_0_11 <= _T_52606[11];
    storeAddrNotKnownFlagsPReg_0_12 <= _T_52606[12];
    storeAddrNotKnownFlagsPReg_0_13 <= _T_52606[13];
    storeAddrNotKnownFlagsPReg_0_14 <= _T_52606[14];
    storeAddrNotKnownFlagsPReg_0_15 <= _T_52606[15];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_53464[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_53464[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_53464[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_53464[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_53464[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_53464[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_53464[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_53464[7];
    storeAddrNotKnownFlagsPReg_1_8 <= _T_53464[8];
    storeAddrNotKnownFlagsPReg_1_9 <= _T_53464[9];
    storeAddrNotKnownFlagsPReg_1_10 <= _T_53464[10];
    storeAddrNotKnownFlagsPReg_1_11 <= _T_53464[11];
    storeAddrNotKnownFlagsPReg_1_12 <= _T_53464[12];
    storeAddrNotKnownFlagsPReg_1_13 <= _T_53464[13];
    storeAddrNotKnownFlagsPReg_1_14 <= _T_53464[14];
    storeAddrNotKnownFlagsPReg_1_15 <= _T_53464[15];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_54322[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_54322[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_54322[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_54322[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_54322[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_54322[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_54322[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_54322[7];
    storeAddrNotKnownFlagsPReg_2_8 <= _T_54322[8];
    storeAddrNotKnownFlagsPReg_2_9 <= _T_54322[9];
    storeAddrNotKnownFlagsPReg_2_10 <= _T_54322[10];
    storeAddrNotKnownFlagsPReg_2_11 <= _T_54322[11];
    storeAddrNotKnownFlagsPReg_2_12 <= _T_54322[12];
    storeAddrNotKnownFlagsPReg_2_13 <= _T_54322[13];
    storeAddrNotKnownFlagsPReg_2_14 <= _T_54322[14];
    storeAddrNotKnownFlagsPReg_2_15 <= _T_54322[15];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_55180[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_55180[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_55180[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_55180[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_55180[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_55180[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_55180[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_55180[7];
    storeAddrNotKnownFlagsPReg_3_8 <= _T_55180[8];
    storeAddrNotKnownFlagsPReg_3_9 <= _T_55180[9];
    storeAddrNotKnownFlagsPReg_3_10 <= _T_55180[10];
    storeAddrNotKnownFlagsPReg_3_11 <= _T_55180[11];
    storeAddrNotKnownFlagsPReg_3_12 <= _T_55180[12];
    storeAddrNotKnownFlagsPReg_3_13 <= _T_55180[13];
    storeAddrNotKnownFlagsPReg_3_14 <= _T_55180[14];
    storeAddrNotKnownFlagsPReg_3_15 <= _T_55180[15];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_56038[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_56038[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_56038[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_56038[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_56038[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_56038[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_56038[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_56038[7];
    storeAddrNotKnownFlagsPReg_4_8 <= _T_56038[8];
    storeAddrNotKnownFlagsPReg_4_9 <= _T_56038[9];
    storeAddrNotKnownFlagsPReg_4_10 <= _T_56038[10];
    storeAddrNotKnownFlagsPReg_4_11 <= _T_56038[11];
    storeAddrNotKnownFlagsPReg_4_12 <= _T_56038[12];
    storeAddrNotKnownFlagsPReg_4_13 <= _T_56038[13];
    storeAddrNotKnownFlagsPReg_4_14 <= _T_56038[14];
    storeAddrNotKnownFlagsPReg_4_15 <= _T_56038[15];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_56896[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_56896[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_56896[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_56896[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_56896[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_56896[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_56896[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_56896[7];
    storeAddrNotKnownFlagsPReg_5_8 <= _T_56896[8];
    storeAddrNotKnownFlagsPReg_5_9 <= _T_56896[9];
    storeAddrNotKnownFlagsPReg_5_10 <= _T_56896[10];
    storeAddrNotKnownFlagsPReg_5_11 <= _T_56896[11];
    storeAddrNotKnownFlagsPReg_5_12 <= _T_56896[12];
    storeAddrNotKnownFlagsPReg_5_13 <= _T_56896[13];
    storeAddrNotKnownFlagsPReg_5_14 <= _T_56896[14];
    storeAddrNotKnownFlagsPReg_5_15 <= _T_56896[15];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_57754[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_57754[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_57754[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_57754[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_57754[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_57754[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_57754[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_57754[7];
    storeAddrNotKnownFlagsPReg_6_8 <= _T_57754[8];
    storeAddrNotKnownFlagsPReg_6_9 <= _T_57754[9];
    storeAddrNotKnownFlagsPReg_6_10 <= _T_57754[10];
    storeAddrNotKnownFlagsPReg_6_11 <= _T_57754[11];
    storeAddrNotKnownFlagsPReg_6_12 <= _T_57754[12];
    storeAddrNotKnownFlagsPReg_6_13 <= _T_57754[13];
    storeAddrNotKnownFlagsPReg_6_14 <= _T_57754[14];
    storeAddrNotKnownFlagsPReg_6_15 <= _T_57754[15];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_58612[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_58612[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_58612[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_58612[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_58612[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_58612[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_58612[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_58612[7];
    storeAddrNotKnownFlagsPReg_7_8 <= _T_58612[8];
    storeAddrNotKnownFlagsPReg_7_9 <= _T_58612[9];
    storeAddrNotKnownFlagsPReg_7_10 <= _T_58612[10];
    storeAddrNotKnownFlagsPReg_7_11 <= _T_58612[11];
    storeAddrNotKnownFlagsPReg_7_12 <= _T_58612[12];
    storeAddrNotKnownFlagsPReg_7_13 <= _T_58612[13];
    storeAddrNotKnownFlagsPReg_7_14 <= _T_58612[14];
    storeAddrNotKnownFlagsPReg_7_15 <= _T_58612[15];
    storeAddrNotKnownFlagsPReg_8_0 <= _T_59470[0];
    storeAddrNotKnownFlagsPReg_8_1 <= _T_59470[1];
    storeAddrNotKnownFlagsPReg_8_2 <= _T_59470[2];
    storeAddrNotKnownFlagsPReg_8_3 <= _T_59470[3];
    storeAddrNotKnownFlagsPReg_8_4 <= _T_59470[4];
    storeAddrNotKnownFlagsPReg_8_5 <= _T_59470[5];
    storeAddrNotKnownFlagsPReg_8_6 <= _T_59470[6];
    storeAddrNotKnownFlagsPReg_8_7 <= _T_59470[7];
    storeAddrNotKnownFlagsPReg_8_8 <= _T_59470[8];
    storeAddrNotKnownFlagsPReg_8_9 <= _T_59470[9];
    storeAddrNotKnownFlagsPReg_8_10 <= _T_59470[10];
    storeAddrNotKnownFlagsPReg_8_11 <= _T_59470[11];
    storeAddrNotKnownFlagsPReg_8_12 <= _T_59470[12];
    storeAddrNotKnownFlagsPReg_8_13 <= _T_59470[13];
    storeAddrNotKnownFlagsPReg_8_14 <= _T_59470[14];
    storeAddrNotKnownFlagsPReg_8_15 <= _T_59470[15];
    storeAddrNotKnownFlagsPReg_9_0 <= _T_60328[0];
    storeAddrNotKnownFlagsPReg_9_1 <= _T_60328[1];
    storeAddrNotKnownFlagsPReg_9_2 <= _T_60328[2];
    storeAddrNotKnownFlagsPReg_9_3 <= _T_60328[3];
    storeAddrNotKnownFlagsPReg_9_4 <= _T_60328[4];
    storeAddrNotKnownFlagsPReg_9_5 <= _T_60328[5];
    storeAddrNotKnownFlagsPReg_9_6 <= _T_60328[6];
    storeAddrNotKnownFlagsPReg_9_7 <= _T_60328[7];
    storeAddrNotKnownFlagsPReg_9_8 <= _T_60328[8];
    storeAddrNotKnownFlagsPReg_9_9 <= _T_60328[9];
    storeAddrNotKnownFlagsPReg_9_10 <= _T_60328[10];
    storeAddrNotKnownFlagsPReg_9_11 <= _T_60328[11];
    storeAddrNotKnownFlagsPReg_9_12 <= _T_60328[12];
    storeAddrNotKnownFlagsPReg_9_13 <= _T_60328[13];
    storeAddrNotKnownFlagsPReg_9_14 <= _T_60328[14];
    storeAddrNotKnownFlagsPReg_9_15 <= _T_60328[15];
    storeAddrNotKnownFlagsPReg_10_0 <= _T_61186[0];
    storeAddrNotKnownFlagsPReg_10_1 <= _T_61186[1];
    storeAddrNotKnownFlagsPReg_10_2 <= _T_61186[2];
    storeAddrNotKnownFlagsPReg_10_3 <= _T_61186[3];
    storeAddrNotKnownFlagsPReg_10_4 <= _T_61186[4];
    storeAddrNotKnownFlagsPReg_10_5 <= _T_61186[5];
    storeAddrNotKnownFlagsPReg_10_6 <= _T_61186[6];
    storeAddrNotKnownFlagsPReg_10_7 <= _T_61186[7];
    storeAddrNotKnownFlagsPReg_10_8 <= _T_61186[8];
    storeAddrNotKnownFlagsPReg_10_9 <= _T_61186[9];
    storeAddrNotKnownFlagsPReg_10_10 <= _T_61186[10];
    storeAddrNotKnownFlagsPReg_10_11 <= _T_61186[11];
    storeAddrNotKnownFlagsPReg_10_12 <= _T_61186[12];
    storeAddrNotKnownFlagsPReg_10_13 <= _T_61186[13];
    storeAddrNotKnownFlagsPReg_10_14 <= _T_61186[14];
    storeAddrNotKnownFlagsPReg_10_15 <= _T_61186[15];
    storeAddrNotKnownFlagsPReg_11_0 <= _T_62044[0];
    storeAddrNotKnownFlagsPReg_11_1 <= _T_62044[1];
    storeAddrNotKnownFlagsPReg_11_2 <= _T_62044[2];
    storeAddrNotKnownFlagsPReg_11_3 <= _T_62044[3];
    storeAddrNotKnownFlagsPReg_11_4 <= _T_62044[4];
    storeAddrNotKnownFlagsPReg_11_5 <= _T_62044[5];
    storeAddrNotKnownFlagsPReg_11_6 <= _T_62044[6];
    storeAddrNotKnownFlagsPReg_11_7 <= _T_62044[7];
    storeAddrNotKnownFlagsPReg_11_8 <= _T_62044[8];
    storeAddrNotKnownFlagsPReg_11_9 <= _T_62044[9];
    storeAddrNotKnownFlagsPReg_11_10 <= _T_62044[10];
    storeAddrNotKnownFlagsPReg_11_11 <= _T_62044[11];
    storeAddrNotKnownFlagsPReg_11_12 <= _T_62044[12];
    storeAddrNotKnownFlagsPReg_11_13 <= _T_62044[13];
    storeAddrNotKnownFlagsPReg_11_14 <= _T_62044[14];
    storeAddrNotKnownFlagsPReg_11_15 <= _T_62044[15];
    storeAddrNotKnownFlagsPReg_12_0 <= _T_62902[0];
    storeAddrNotKnownFlagsPReg_12_1 <= _T_62902[1];
    storeAddrNotKnownFlagsPReg_12_2 <= _T_62902[2];
    storeAddrNotKnownFlagsPReg_12_3 <= _T_62902[3];
    storeAddrNotKnownFlagsPReg_12_4 <= _T_62902[4];
    storeAddrNotKnownFlagsPReg_12_5 <= _T_62902[5];
    storeAddrNotKnownFlagsPReg_12_6 <= _T_62902[6];
    storeAddrNotKnownFlagsPReg_12_7 <= _T_62902[7];
    storeAddrNotKnownFlagsPReg_12_8 <= _T_62902[8];
    storeAddrNotKnownFlagsPReg_12_9 <= _T_62902[9];
    storeAddrNotKnownFlagsPReg_12_10 <= _T_62902[10];
    storeAddrNotKnownFlagsPReg_12_11 <= _T_62902[11];
    storeAddrNotKnownFlagsPReg_12_12 <= _T_62902[12];
    storeAddrNotKnownFlagsPReg_12_13 <= _T_62902[13];
    storeAddrNotKnownFlagsPReg_12_14 <= _T_62902[14];
    storeAddrNotKnownFlagsPReg_12_15 <= _T_62902[15];
    storeAddrNotKnownFlagsPReg_13_0 <= _T_63760[0];
    storeAddrNotKnownFlagsPReg_13_1 <= _T_63760[1];
    storeAddrNotKnownFlagsPReg_13_2 <= _T_63760[2];
    storeAddrNotKnownFlagsPReg_13_3 <= _T_63760[3];
    storeAddrNotKnownFlagsPReg_13_4 <= _T_63760[4];
    storeAddrNotKnownFlagsPReg_13_5 <= _T_63760[5];
    storeAddrNotKnownFlagsPReg_13_6 <= _T_63760[6];
    storeAddrNotKnownFlagsPReg_13_7 <= _T_63760[7];
    storeAddrNotKnownFlagsPReg_13_8 <= _T_63760[8];
    storeAddrNotKnownFlagsPReg_13_9 <= _T_63760[9];
    storeAddrNotKnownFlagsPReg_13_10 <= _T_63760[10];
    storeAddrNotKnownFlagsPReg_13_11 <= _T_63760[11];
    storeAddrNotKnownFlagsPReg_13_12 <= _T_63760[12];
    storeAddrNotKnownFlagsPReg_13_13 <= _T_63760[13];
    storeAddrNotKnownFlagsPReg_13_14 <= _T_63760[14];
    storeAddrNotKnownFlagsPReg_13_15 <= _T_63760[15];
    storeAddrNotKnownFlagsPReg_14_0 <= _T_64618[0];
    storeAddrNotKnownFlagsPReg_14_1 <= _T_64618[1];
    storeAddrNotKnownFlagsPReg_14_2 <= _T_64618[2];
    storeAddrNotKnownFlagsPReg_14_3 <= _T_64618[3];
    storeAddrNotKnownFlagsPReg_14_4 <= _T_64618[4];
    storeAddrNotKnownFlagsPReg_14_5 <= _T_64618[5];
    storeAddrNotKnownFlagsPReg_14_6 <= _T_64618[6];
    storeAddrNotKnownFlagsPReg_14_7 <= _T_64618[7];
    storeAddrNotKnownFlagsPReg_14_8 <= _T_64618[8];
    storeAddrNotKnownFlagsPReg_14_9 <= _T_64618[9];
    storeAddrNotKnownFlagsPReg_14_10 <= _T_64618[10];
    storeAddrNotKnownFlagsPReg_14_11 <= _T_64618[11];
    storeAddrNotKnownFlagsPReg_14_12 <= _T_64618[12];
    storeAddrNotKnownFlagsPReg_14_13 <= _T_64618[13];
    storeAddrNotKnownFlagsPReg_14_14 <= _T_64618[14];
    storeAddrNotKnownFlagsPReg_14_15 <= _T_64618[15];
    storeAddrNotKnownFlagsPReg_15_0 <= _T_65476[0];
    storeAddrNotKnownFlagsPReg_15_1 <= _T_65476[1];
    storeAddrNotKnownFlagsPReg_15_2 <= _T_65476[2];
    storeAddrNotKnownFlagsPReg_15_3 <= _T_65476[3];
    storeAddrNotKnownFlagsPReg_15_4 <= _T_65476[4];
    storeAddrNotKnownFlagsPReg_15_5 <= _T_65476[5];
    storeAddrNotKnownFlagsPReg_15_6 <= _T_65476[6];
    storeAddrNotKnownFlagsPReg_15_7 <= _T_65476[7];
    storeAddrNotKnownFlagsPReg_15_8 <= _T_65476[8];
    storeAddrNotKnownFlagsPReg_15_9 <= _T_65476[9];
    storeAddrNotKnownFlagsPReg_15_10 <= _T_65476[10];
    storeAddrNotKnownFlagsPReg_15_11 <= _T_65476[11];
    storeAddrNotKnownFlagsPReg_15_12 <= _T_65476[12];
    storeAddrNotKnownFlagsPReg_15_13 <= _T_65476[13];
    storeAddrNotKnownFlagsPReg_15_14 <= _T_65476[14];
    storeAddrNotKnownFlagsPReg_15_15 <= _T_65476[15];
    shiftedStoreDataKnownPReg_0 <= _T_5972[0];
    shiftedStoreDataKnownPReg_1 <= _T_5972[1];
    shiftedStoreDataKnownPReg_2 <= _T_5972[2];
    shiftedStoreDataKnownPReg_3 <= _T_5972[3];
    shiftedStoreDataKnownPReg_4 <= _T_5972[4];
    shiftedStoreDataKnownPReg_5 <= _T_5972[5];
    shiftedStoreDataKnownPReg_6 <= _T_5972[6];
    shiftedStoreDataKnownPReg_7 <= _T_5972[7];
    shiftedStoreDataKnownPReg_8 <= _T_5972[8];
    shiftedStoreDataKnownPReg_9 <= _T_5972[9];
    shiftedStoreDataKnownPReg_10 <= _T_5972[10];
    shiftedStoreDataKnownPReg_11 <= _T_5972[11];
    shiftedStoreDataKnownPReg_12 <= _T_5972[12];
    shiftedStoreDataKnownPReg_13 <= _T_5972[13];
    shiftedStoreDataKnownPReg_14 <= _T_5972[14];
    shiftedStoreDataKnownPReg_15 <= _T_5972[15];
    shiftedStoreDataQPreg_0 <= _T_5115[31:0];
    shiftedStoreDataQPreg_1 <= _T_5115[63:32];
    shiftedStoreDataQPreg_2 <= _T_5115[95:64];
    shiftedStoreDataQPreg_3 <= _T_5115[127:96];
    shiftedStoreDataQPreg_4 <= _T_5115[159:128];
    shiftedStoreDataQPreg_5 <= _T_5115[191:160];
    shiftedStoreDataQPreg_6 <= _T_5115[223:192];
    shiftedStoreDataQPreg_7 <= _T_5115[255:224];
    shiftedStoreDataQPreg_8 <= _T_5115[287:256];
    shiftedStoreDataQPreg_9 <= _T_5115[319:288];
    shiftedStoreDataQPreg_10 <= _T_5115[351:320];
    shiftedStoreDataQPreg_11 <= _T_5115[383:352];
    shiftedStoreDataQPreg_12 <= _T_5115[415:384];
    shiftedStoreDataQPreg_13 <= _T_5115[447:416];
    shiftedStoreDataQPreg_14 <= _T_5115[479:448];
    shiftedStoreDataQPreg_15 <= _T_5115[511:480];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    addrKnownPReg_8 <= addrKnown_8;
    addrKnownPReg_9 <= addrKnown_9;
    addrKnownPReg_10 <= addrKnown_10;
    addrKnownPReg_11 <= addrKnown_11;
    addrKnownPReg_12 <= addrKnown_12;
    addrKnownPReg_13 <= addrKnown_13;
    addrKnownPReg_14 <= addrKnown_14;
    addrKnownPReg_15 <= addrKnown_15;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    dataKnownPReg_8 <= dataKnown_8;
    dataKnownPReg_9 <= dataKnown_9;
    dataKnownPReg_10 <= dataKnown_10;
    dataKnownPReg_11 <= dataKnown_11;
    dataKnownPReg_12 <= dataKnown_12;
    dataKnownPReg_13 <= dataKnown_13;
    dataKnownPReg_14 <= dataKnown_14;
    dataKnownPReg_15 <= dataKnown_15;
    if (reset) begin
      prevPriorityRequest_15 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_15 <= priorityLoadRequest_15;
      end else begin
        prevPriorityRequest_15 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_14 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_14 <= priorityLoadRequest_14;
      end else begin
        prevPriorityRequest_14 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_13 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_13 <= priorityLoadRequest_13;
      end else begin
        prevPriorityRequest_13 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_12 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_12 <= priorityLoadRequest_12;
      end else begin
        prevPriorityRequest_12 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_11 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_11 <= priorityLoadRequest_11;
      end else begin
        prevPriorityRequest_11 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_10 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_10 <= priorityLoadRequest_10;
      end else begin
        prevPriorityRequest_10 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_9 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_9 <= priorityLoadRequest_9;
      end else begin
        prevPriorityRequest_9 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_8 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_8 <= priorityLoadRequest_8;
      end else begin
        prevPriorityRequest_8 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_7 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_7 <= priorityLoadRequest_7;
      end else begin
        prevPriorityRequest_7 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_6 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_6 <= priorityLoadRequest_6;
      end else begin
        prevPriorityRequest_6 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_5 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_5 <= priorityLoadRequest_5;
      end else begin
        prevPriorityRequest_5 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_4 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_4 <= priorityLoadRequest_4;
      end else begin
        prevPriorityRequest_4 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_3 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_3 <= priorityLoadRequest_3;
      end else begin
        prevPriorityRequest_3 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_2 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_2 <= priorityLoadRequest_2;
      end else begin
        prevPriorityRequest_2 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_1 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_1 <= priorityLoadRequest_1;
      end else begin
        prevPriorityRequest_1 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_0 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_0 <= priorityLoadRequest_0;
      end else begin
        prevPriorityRequest_0 <= 1'h0;
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_E( // @[:@45077.2]
  output [3:0] io_bbLoadOffsets_0, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_1, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_2, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_3, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_4, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_5, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_6, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_7, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_8, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_9, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_10, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_11, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_12, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_13, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_14, // @[:@45080.4]
  output [3:0] io_bbLoadOffsets_15, // @[:@45080.4]
  output       io_bbNumLoads, // @[:@45080.4]
  input  [3:0] io_loadTail, // @[:@45080.4]
  input  [3:0] io_loadHead, // @[:@45080.4]
  input        io_loadEmpty, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_0, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_1, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_2, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_3, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_4, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_5, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_6, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_7, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_8, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_9, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_10, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_11, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_12, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_13, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_14, // @[:@45080.4]
  output [3:0] io_bbStoreOffsets_15, // @[:@45080.4]
  output       io_bbStorePorts_0, // @[:@45080.4]
  output [1:0] io_bbNumStores, // @[:@45080.4]
  input  [3:0] io_storeTail, // @[:@45080.4]
  input  [3:0] io_storeHead, // @[:@45080.4]
  input        io_storeEmpty, // @[:@45080.4]
  output       io_bbStart, // @[:@45080.4]
  input        io_bbStartSignals_0, // @[:@45080.4]
  input        io_bbStartSignals_1, // @[:@45080.4]
  output       io_readyToPrevious_0, // @[:@45080.4]
  output       io_readyToPrevious_1, // @[:@45080.4]
  output       io_loadPortsEnable_0, // @[:@45080.4]
  output       io_storePortsEnable_0, // @[:@45080.4]
  output       io_storePortsEnable_1 // @[:@45080.4]
);
  wire  _T_246; // @[GroupAllocator.scala 42:25:@45083.4]
  wire  _T_247; // @[GroupAllocator.scala 42:16:@45084.4]
  wire [4:0] _GEN_68; // @[GroupAllocator.scala 43:36:@45086.6]
  wire [5:0] _T_249; // @[GroupAllocator.scala 43:36:@45086.6]
  wire [5:0] _T_250; // @[GroupAllocator.scala 43:36:@45087.6]
  wire [4:0] _T_251; // @[GroupAllocator.scala 43:36:@45088.6]
  wire [4:0] _GEN_69; // @[GroupAllocator.scala 43:43:@45089.6]
  wire [5:0] _T_252; // @[GroupAllocator.scala 43:43:@45089.6]
  wire [4:0] _T_253; // @[GroupAllocator.scala 43:43:@45090.6]
  wire [4:0] _T_254; // @[GroupAllocator.scala 45:22:@45094.6]
  wire [4:0] _T_255; // @[GroupAllocator.scala 45:22:@45095.6]
  wire [3:0] _T_256; // @[GroupAllocator.scala 45:22:@45096.6]
  wire [4:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@45085.4]
  wire  _T_258; // @[GroupAllocator.scala 42:25:@45100.4]
  wire  _T_259; // @[GroupAllocator.scala 42:16:@45101.4]
  wire [4:0] _GEN_70; // @[GroupAllocator.scala 43:36:@45103.6]
  wire [5:0] _T_261; // @[GroupAllocator.scala 43:36:@45103.6]
  wire [5:0] _T_262; // @[GroupAllocator.scala 43:36:@45104.6]
  wire [4:0] _T_263; // @[GroupAllocator.scala 43:36:@45105.6]
  wire [4:0] _GEN_71; // @[GroupAllocator.scala 43:43:@45106.6]
  wire [5:0] _T_264; // @[GroupAllocator.scala 43:43:@45106.6]
  wire [4:0] _T_265; // @[GroupAllocator.scala 43:43:@45107.6]
  wire [4:0] _T_266; // @[GroupAllocator.scala 45:22:@45111.6]
  wire [4:0] _T_267; // @[GroupAllocator.scala 45:22:@45112.6]
  wire [3:0] _T_268; // @[GroupAllocator.scala 45:22:@45113.6]
  wire [4:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@45102.4]
  wire  _T_270; // @[GroupAllocator.scala 54:19:@45116.4]
  wire  _T_277; // @[GroupAllocator.scala 54:50:@45120.4]
  wire  possibleAllocations_0; // @[GroupAllocator.scala 56:106:@45127.4]
  wire  possibleAllocations_1; // @[GroupAllocator.scala 56:106:@45128.4]
  wire  allocatedBBIdx; // @[Mux.scala 31:69:@45132.4]
  wire  _T_305; // @[GroupAllocator.scala 78:44:@45139.4]
  wire  _T_472; // @[Mux.scala 46:16:@45283.6]
  wire  _T_481; // @[Mux.scala 46:16:@45288.6]
  wire [5:0] _T_903; // @[GroupAllocator.scala 110:34:@45449.6]
  wire [4:0] _T_904; // @[GroupAllocator.scala 110:34:@45450.6]
  wire [5:0] _T_906; // @[GroupAllocator.scala 110:55:@45451.6]
  wire [5:0] _T_907; // @[GroupAllocator.scala 110:55:@45452.6]
  wire [4:0] _T_908; // @[GroupAllocator.scala 110:55:@45453.6]
  wire [5:0] _T_910; // @[util.scala 10:8:@45454.6]
  wire [5:0] _GEN_0; // @[util.scala 10:14:@45455.6]
  wire [4:0] _T_911; // @[util.scala 10:14:@45455.6]
  wire [3:0] _T_1161; // @[GroupAllocator.scala 110:90:@45617.6 GroupAllocator.scala 110:90:@45618.6]
  wire [3:0] _T_1395_0; // @[Mux.scala 46:16:@45772.6]
  wire [3:0] _T_1432_0; // @[Mux.scala 46:16:@45774.6]
  wire [5:0] _T_1509; // @[GroupAllocator.scala 115:33:@45808.6]
  wire [4:0] _T_1510; // @[GroupAllocator.scala 115:33:@45809.6]
  wire [5:0] _T_1512; // @[GroupAllocator.scala 115:54:@45810.6]
  wire [5:0] _T_1513; // @[GroupAllocator.scala 115:54:@45811.6]
  wire [4:0] _T_1514; // @[GroupAllocator.scala 115:54:@45812.6]
  wire [5:0] _T_1516; // @[util.scala 10:8:@45813.6]
  wire [5:0] _GEN_1; // @[util.scala 10:14:@45814.6]
  wire [4:0] _T_1517; // @[util.scala 10:14:@45814.6]
  wire [5:0] _T_1763; // @[util.scala 10:8:@45974.6]
  wire [5:0] _GEN_2; // @[util.scala 10:14:@45975.6]
  wire [4:0] _T_1764; // @[util.scala 10:14:@45975.6]
  wire [3:0] _T_1767; // @[GroupAllocator.scala 115:89:@45976.6 GroupAllocator.scala 115:89:@45977.6]
  wire [3:0] _T_2001_0; // @[Mux.scala 46:16:@46131.6]
  wire [3:0] _T_1781; // @[GroupAllocator.scala 115:89:@45985.6 GroupAllocator.scala 115:89:@45986.6]
  wire [3:0] _T_2001_1; // @[Mux.scala 46:16:@46131.6]
  wire [3:0] _T_2038_0; // @[Mux.scala 46:16:@46133.6]
  wire [3:0] _T_2038_1; // @[Mux.scala 46:16:@46133.6]
  assign _T_246 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@45083.4]
  assign _T_247 = io_loadEmpty | _T_246; // @[GroupAllocator.scala 42:16:@45084.4]
  assign _GEN_68 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@45086.6]
  assign _T_249 = 5'h10 - _GEN_68; // @[GroupAllocator.scala 43:36:@45086.6]
  assign _T_250 = $unsigned(_T_249); // @[GroupAllocator.scala 43:36:@45087.6]
  assign _T_251 = _T_250[4:0]; // @[GroupAllocator.scala 43:36:@45088.6]
  assign _GEN_69 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@45089.6]
  assign _T_252 = _T_251 + _GEN_69; // @[GroupAllocator.scala 43:43:@45089.6]
  assign _T_253 = _T_251 + _GEN_69; // @[GroupAllocator.scala 43:43:@45090.6]
  assign _T_254 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@45094.6]
  assign _T_255 = $unsigned(_T_254); // @[GroupAllocator.scala 45:22:@45095.6]
  assign _T_256 = _T_255[3:0]; // @[GroupAllocator.scala 45:22:@45096.6]
  assign emptyLoadSlots = _T_247 ? _T_253 : {{1'd0}, _T_256}; // @[GroupAllocator.scala 42:34:@45085.4]
  assign _T_258 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@45100.4]
  assign _T_259 = io_storeEmpty | _T_258; // @[GroupAllocator.scala 42:16:@45101.4]
  assign _GEN_70 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@45103.6]
  assign _T_261 = 5'h10 - _GEN_70; // @[GroupAllocator.scala 43:36:@45103.6]
  assign _T_262 = $unsigned(_T_261); // @[GroupAllocator.scala 43:36:@45104.6]
  assign _T_263 = _T_262[4:0]; // @[GroupAllocator.scala 43:36:@45105.6]
  assign _GEN_71 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@45106.6]
  assign _T_264 = _T_263 + _GEN_71; // @[GroupAllocator.scala 43:43:@45106.6]
  assign _T_265 = _T_263 + _GEN_71; // @[GroupAllocator.scala 43:43:@45107.6]
  assign _T_266 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@45111.6]
  assign _T_267 = $unsigned(_T_266); // @[GroupAllocator.scala 45:22:@45112.6]
  assign _T_268 = _T_267[3:0]; // @[GroupAllocator.scala 45:22:@45113.6]
  assign emptyStoreSlots = _T_259 ? _T_265 : {{1'd0}, _T_268}; // @[GroupAllocator.scala 42:34:@45102.4]
  assign _T_270 = 5'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 54:19:@45116.4]
  assign _T_277 = 5'h1 <= emptyLoadSlots; // @[GroupAllocator.scala 54:50:@45120.4]
  assign possibleAllocations_0 = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 56:106:@45127.4]
  assign possibleAllocations_1 = io_readyToPrevious_1 & io_bbStartSignals_1; // @[GroupAllocator.scala 56:106:@45128.4]
  assign allocatedBBIdx = possibleAllocations_0 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@45132.4]
  assign _T_305 = 1'h0 == allocatedBBIdx; // @[GroupAllocator.scala 78:44:@45139.4]
  assign _T_472 = _T_305 ? 1'h0 : allocatedBBIdx; // @[Mux.scala 46:16:@45283.6]
  assign _T_481 = _T_305 ? 1'h1 : allocatedBBIdx; // @[Mux.scala 46:16:@45288.6]
  assign _T_903 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@45449.6]
  assign _T_904 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@45450.6]
  assign _T_906 = _T_904 - 5'h1; // @[GroupAllocator.scala 110:55:@45451.6]
  assign _T_907 = $unsigned(_T_906); // @[GroupAllocator.scala 110:55:@45452.6]
  assign _T_908 = _T_907[4:0]; // @[GroupAllocator.scala 110:55:@45453.6]
  assign _T_910 = {{1'd0}, _T_908}; // @[util.scala 10:8:@45454.6]
  assign _GEN_0 = _T_910 % 6'h10; // @[util.scala 10:14:@45455.6]
  assign _T_911 = _GEN_0[4:0]; // @[util.scala 10:14:@45455.6]
  assign _T_1161 = _T_911[3:0]; // @[GroupAllocator.scala 110:90:@45617.6 GroupAllocator.scala 110:90:@45618.6]
  assign _T_1395_0 = allocatedBBIdx ? _T_1161 : 4'h0; // @[Mux.scala 46:16:@45772.6]
  assign _T_1432_0 = _T_305 ? _T_1161 : _T_1395_0; // @[Mux.scala 46:16:@45774.6]
  assign _T_1509 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@45808.6]
  assign _T_1510 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@45809.6]
  assign _T_1512 = _T_1510 - 5'h1; // @[GroupAllocator.scala 115:54:@45810.6]
  assign _T_1513 = $unsigned(_T_1512); // @[GroupAllocator.scala 115:54:@45811.6]
  assign _T_1514 = _T_1513[4:0]; // @[GroupAllocator.scala 115:54:@45812.6]
  assign _T_1516 = {{1'd0}, _T_1514}; // @[util.scala 10:8:@45813.6]
  assign _GEN_1 = _T_1516 % 6'h10; // @[util.scala 10:14:@45814.6]
  assign _T_1517 = _GEN_1[4:0]; // @[util.scala 10:14:@45814.6]
  assign _T_1763 = 5'h1 + _T_1514; // @[util.scala 10:8:@45974.6]
  assign _GEN_2 = _T_1763 % 6'h10; // @[util.scala 10:14:@45975.6]
  assign _T_1764 = _GEN_2[4:0]; // @[util.scala 10:14:@45975.6]
  assign _T_1767 = _T_1764[3:0]; // @[GroupAllocator.scala 115:89:@45976.6 GroupAllocator.scala 115:89:@45977.6]
  assign _T_2001_0 = allocatedBBIdx ? _T_1767 : 4'h0; // @[Mux.scala 46:16:@46131.6]
  assign _T_1781 = _T_1517[3:0]; // @[GroupAllocator.scala 115:89:@45985.6 GroupAllocator.scala 115:89:@45986.6]
  assign _T_2001_1 = allocatedBBIdx ? _T_1781 : 4'h0; // @[Mux.scala 46:16:@46131.6]
  assign _T_2038_0 = _T_305 ? _T_1781 : _T_2001_0; // @[Mux.scala 46:16:@46133.6]
  assign _T_2038_1 = _T_305 ? _T_1781 : _T_2001_1; // @[Mux.scala 46:16:@46133.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45230.4 GroupAllocator.scala 106:22:@45775.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45231.4 GroupAllocator.scala 106:22:@45776.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45232.4 GroupAllocator.scala 106:22:@45777.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45233.4 GroupAllocator.scala 106:22:@45778.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45234.4 GroupAllocator.scala 106:22:@45779.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45235.4 GroupAllocator.scala 106:22:@45780.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45236.4 GroupAllocator.scala 106:22:@45781.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45237.4 GroupAllocator.scala 106:22:@45782.6]
  assign io_bbLoadOffsets_8 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45238.4 GroupAllocator.scala 106:22:@45783.6]
  assign io_bbLoadOffsets_9 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45239.4 GroupAllocator.scala 106:22:@45784.6]
  assign io_bbLoadOffsets_10 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45240.4 GroupAllocator.scala 106:22:@45785.6]
  assign io_bbLoadOffsets_11 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45241.4 GroupAllocator.scala 106:22:@45786.6]
  assign io_bbLoadOffsets_12 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45242.4 GroupAllocator.scala 106:22:@45787.6]
  assign io_bbLoadOffsets_13 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45243.4 GroupAllocator.scala 106:22:@45788.6]
  assign io_bbLoadOffsets_14 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45244.4 GroupAllocator.scala 106:22:@45789.6]
  assign io_bbLoadOffsets_15 = io_bbStart ? _T_1432_0 : 4'h0; // @[GroupAllocator.scala 89:20:@45245.4 GroupAllocator.scala 106:22:@45790.6]
  assign io_bbNumLoads = io_bbStart ? _T_472 : 1'h0; // @[GroupAllocator.scala 85:17:@45145.4 GroupAllocator.scala 93:19:@45284.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_2038_0 : 4'h0; // @[GroupAllocator.scala 90:21:@45263.4 GroupAllocator.scala 111:23:@46134.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45264.4 GroupAllocator.scala 111:23:@46135.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45265.4 GroupAllocator.scala 111:23:@46136.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45266.4 GroupAllocator.scala 111:23:@46137.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45267.4 GroupAllocator.scala 111:23:@46138.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45268.4 GroupAllocator.scala 111:23:@46139.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45269.4 GroupAllocator.scala 111:23:@46140.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45270.4 GroupAllocator.scala 111:23:@46141.6]
  assign io_bbStoreOffsets_8 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45271.4 GroupAllocator.scala 111:23:@46142.6]
  assign io_bbStoreOffsets_9 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45272.4 GroupAllocator.scala 111:23:@46143.6]
  assign io_bbStoreOffsets_10 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45273.4 GroupAllocator.scala 111:23:@46144.6]
  assign io_bbStoreOffsets_11 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45274.4 GroupAllocator.scala 111:23:@46145.6]
  assign io_bbStoreOffsets_12 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45275.4 GroupAllocator.scala 111:23:@46146.6]
  assign io_bbStoreOffsets_13 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45276.4 GroupAllocator.scala 111:23:@46147.6]
  assign io_bbStoreOffsets_14 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45277.4 GroupAllocator.scala 111:23:@46148.6]
  assign io_bbStoreOffsets_15 = io_bbStart ? _T_2038_1 : 4'h0; // @[GroupAllocator.scala 90:21:@45278.4 GroupAllocator.scala 111:23:@46149.6]
  assign io_bbStorePorts_0 = io_bbStart ? _T_472 : 1'h0; // @[GroupAllocator.scala 88:19:@45197.4 GroupAllocator.scala 100:21:@45416.6]
  assign io_bbNumStores = io_bbStart ? {{1'd0}, _T_481} : 2'h0; // @[GroupAllocator.scala 86:18:@45146.4 GroupAllocator.scala 94:20:@45289.6]
  assign io_bbStart = possibleAllocations_0 | possibleAllocations_1; // @[GroupAllocator.scala 59:14:@45135.4]
  assign io_readyToPrevious_0 = 5'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 53:22:@45125.4]
  assign io_readyToPrevious_1 = _T_270 & _T_277; // @[GroupAllocator.scala 53:22:@45126.4]
  assign io_loadPortsEnable_0 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 69:29:@45138.4]
  assign io_storePortsEnable_0 = _T_305 & io_bbStart; // @[GroupAllocator.scala 78:30:@45141.4]
  assign io_storePortsEnable_1 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 78:30:@45144.4]
endmodule
module LOAD_PORT_LSQ_E( // @[:@46152.2]
  input         clock, // @[:@46153.4]
  input         reset, // @[:@46154.4]
  output        io_addrFromPrev_ready, // @[:@46155.4]
  input         io_addrFromPrev_valid, // @[:@46155.4]
  input  [31:0] io_addrFromPrev_bits, // @[:@46155.4]
  input         io_portEnable, // @[:@46155.4]
  input         io_dataToNext_ready, // @[:@46155.4]
  output        io_dataToNext_valid, // @[:@46155.4]
  output [31:0] io_dataToNext_bits, // @[:@46155.4]
  output        io_loadAddrEnable, // @[:@46155.4]
  output [31:0] io_addrToLoadQueue, // @[:@46155.4]
  output        io_dataFromLoadQueue_ready, // @[:@46155.4]
  input         io_dataFromLoadQueue_valid, // @[:@46155.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@46155.4]
);
  reg [4:0] cnt; // @[LoadPort.scala 23:20:@46157.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@46158.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@46159.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@46160.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@46161.4]
  wire [5:0] _T_50; // @[LoadPort.scala 27:16:@46163.6]
  wire [4:0] _T_51; // @[LoadPort.scala 27:16:@46164.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@46168.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@46169.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@46170.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@46171.6]
  wire [5:0] _T_59; // @[LoadPort.scala 29:16:@46173.8]
  wire [5:0] _T_60; // @[LoadPort.scala 29:16:@46174.8]
  wire [4:0] _T_61; // @[LoadPort.scala 29:16:@46175.8]
  wire [4:0] _GEN_0; // @[LoadPort.scala 28:66:@46172.6]
  wire [4:0] _GEN_1; // @[LoadPort.scala 26:75:@46162.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@46179.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@46158.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@46159.4]
  assign _T_47 = cnt != 5'h10; // @[LoadPort.scala 26:51:@46160.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@46161.4]
  assign _T_50 = cnt + 5'h1; // @[LoadPort.scala 27:16:@46163.6]
  assign _T_51 = cnt + 5'h1; // @[LoadPort.scala 27:16:@46164.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@46168.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@46169.6]
  assign _T_56 = cnt != 5'h0; // @[LoadPort.scala 28:57:@46170.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@46171.6]
  assign _T_59 = cnt - 5'h1; // @[LoadPort.scala 29:16:@46173.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@46174.8]
  assign _T_61 = _T_60[4:0]; // @[LoadPort.scala 29:16:@46175.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@46172.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@46162.4]
  assign _T_63 = cnt > 5'h0; // @[LoadPort.scala 33:28:@46179.4]
  assign io_addrFromPrev_ready = cnt > 5'h0; // @[LoadPort.scala 34:25:@46183.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@46185.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@46184.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@46181.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@46178.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@46186.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_E( // @[:@46188.2]
  input         clock, // @[:@46189.4]
  input         reset, // @[:@46190.4]
  output        io_dataFromPrev_ready, // @[:@46191.4]
  input         io_dataFromPrev_valid, // @[:@46191.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@46191.4]
  input         io_portEnable, // @[:@46191.4]
  output        io_storeDataEnable, // @[:@46191.4]
  output [31:0] io_dataToStoreQueue // @[:@46191.4]
);
  reg [4:0] cnt; // @[StoreDataPort.scala 21:20:@46193.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@46194.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@46195.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@46196.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@46197.4]
  wire [5:0] _T_32; // @[StoreDataPort.scala 25:16:@46199.6]
  wire [4:0] _T_33; // @[StoreDataPort.scala 25:16:@46200.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@46204.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@46205.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@46206.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@46207.6]
  wire [5:0] _T_41; // @[StoreDataPort.scala 27:16:@46209.8]
  wire [5:0] _T_42; // @[StoreDataPort.scala 27:16:@46210.8]
  wire [4:0] _T_43; // @[StoreDataPort.scala 27:16:@46211.8]
  wire [4:0] _GEN_0; // @[StoreDataPort.scala 26:67:@46208.6]
  wire [4:0] _GEN_1; // @[StoreDataPort.scala 24:76:@46198.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@46215.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@46194.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@46195.4]
  assign _T_29 = cnt != 5'h10; // @[StoreDataPort.scala 24:52:@46196.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@46197.4]
  assign _T_32 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@46199.6]
  assign _T_33 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@46200.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@46204.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@46205.6]
  assign _T_38 = cnt != 5'h0; // @[StoreDataPort.scala 26:58:@46206.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@46207.6]
  assign _T_41 = cnt - 5'h1; // @[StoreDataPort.scala 27:16:@46209.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@46210.8]
  assign _T_43 = _T_42[4:0]; // @[StoreDataPort.scala 27:16:@46211.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@46208.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@46198.4]
  assign _T_45 = cnt > 5'h0; // @[StoreDataPort.scala 31:29:@46215.4]
  assign io_dataFromPrev_ready = cnt > 5'h0; // @[StoreDataPort.scala 32:25:@46219.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@46217.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@46214.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_E( // @[:@46320.2]
  input         clock, // @[:@46321.4]
  input         reset, // @[:@46322.4]
  output [31:0] io_storeDataOut, // @[:@46323.4]
  output [31:0] io_storeAddrOut, // @[:@46323.4]
  output        io_storeEnable, // @[:@46323.4]
  input         io_memIsReadyForStores, // @[:@46323.4]
  input  [31:0] io_loadDataIn, // @[:@46323.4]
  output [31:0] io_loadAddrOut, // @[:@46323.4]
  output        io_loadEnable, // @[:@46323.4]
  input         io_memIsReadyForLoads, // @[:@46323.4]
  input         io_bbpValids_0, // @[:@46323.4]
  input         io_bbpValids_1, // @[:@46323.4]
  output        io_bbReadyToPrevs_0, // @[:@46323.4]
  output        io_bbReadyToPrevs_1, // @[:@46323.4]
  output        io_rdPortsPrev_0_ready, // @[:@46323.4]
  input         io_rdPortsPrev_0_valid, // @[:@46323.4]
  input  [31:0] io_rdPortsPrev_0_bits, // @[:@46323.4]
  input         io_rdPortsNext_0_ready, // @[:@46323.4]
  output        io_rdPortsNext_0_valid, // @[:@46323.4]
  output [31:0] io_rdPortsNext_0_bits, // @[:@46323.4]
  output        io_wrAddrPorts_0_ready, // @[:@46323.4]
  input         io_wrAddrPorts_0_valid, // @[:@46323.4]
  input  [31:0] io_wrAddrPorts_0_bits, // @[:@46323.4]
  output        io_wrAddrPorts_1_ready, // @[:@46323.4]
  input         io_wrAddrPorts_1_valid, // @[:@46323.4]
  input  [31:0] io_wrAddrPorts_1_bits, // @[:@46323.4]
  output        io_wrDataPorts_0_ready, // @[:@46323.4]
  input         io_wrDataPorts_0_valid, // @[:@46323.4]
  input  [31:0] io_wrDataPorts_0_bits, // @[:@46323.4]
  output        io_wrDataPorts_1_ready, // @[:@46323.4]
  input         io_wrDataPorts_1_valid, // @[:@46323.4]
  input  [31:0] io_wrDataPorts_1_bits, // @[:@46323.4]
  output        io_Empty_Valid // @[:@46323.4]
);
  wire  storeQ_clock; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_reset; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_bbStart; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_bbStoreOffsets_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_bbStorePorts_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_bbNumStores; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_storeTail; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_storeHead; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeEmpty; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_loadTail; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [3:0] storeQ_io_loadHead; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadEmpty; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadAddressDone_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_loadDataDone_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_loadAddressQueue_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeDataEnable_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_dataFromStorePorts_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeAddrEnable_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_addressFromStorePorts_0; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_addressFromStorePorts_1; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 72:22:@46354.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  storeQ_io_memIsReadyForStores; // @[LSQBRAM.scala 72:22:@46354.4]
  wire  loadQ_clock; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_reset; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_bbStart; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_bbLoadOffsets_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_bbNumLoads; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_loadTail; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_loadHead; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadEmpty; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_storeTail; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] loadQ_io_storeHead; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeEmpty; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeAddrDone_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_storeDataDone_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_storeDataQueue_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_0; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [31:0] loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 73:21:@46357.4]
  wire  loadQ_io_memIsReadyForLoads; // @[LSQBRAM.scala 73:21:@46357.4]
  wire [3:0] GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_bbNumLoads; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_loadTail; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_loadHead; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_loadEmpty; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_bbStorePorts_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [1:0] GA_io_bbNumStores; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_storeTail; // @[LSQBRAM.scala 74:18:@46360.4]
  wire [3:0] GA_io_storeHead; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_storeEmpty; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_bbStart; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_bbStartSignals_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_bbStartSignals_1; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_readyToPrevious_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_readyToPrevious_1; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_storePortsEnable_0; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  GA_io_storePortsEnable_1; // @[LSQBRAM.scala 74:18:@46360.4]
  wire  LOAD_PORT_LSQ_E_clock; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_reset; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@46363.4]
  wire [31:0] LOAD_PORT_LSQ_E_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_portEnable; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@46363.4]
  wire [31:0] LOAD_PORT_LSQ_E_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@46363.4]
  wire [31:0] LOAD_PORT_LSQ_E_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  LOAD_PORT_LSQ_E_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@46363.4]
  wire [31:0] LOAD_PORT_LSQ_E_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@46363.4]
  wire  STORE_DATA_PORT_LSQ_E_clock; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_reset; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@46379.4]
  wire [31:0] STORE_DATA_PORT_LSQ_E_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_io_portEnable; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@46379.4]
  wire [31:0] STORE_DATA_PORT_LSQ_E_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@46379.4]
  wire  STORE_DATA_PORT_LSQ_E_1_clock; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_DATA_PORT_LSQ_E_1_reset; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@46382.4]
  wire [31:0] STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_DATA_PORT_LSQ_E_1_io_portEnable; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_DATA_PORT_LSQ_E_1_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@46382.4]
  wire [31:0] STORE_DATA_PORT_LSQ_E_1_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@46382.4]
  wire  STORE_ADDR_PORT_LSQ_E_clock; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_reset; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@46398.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_io_portEnable; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@46398.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_E_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@46398.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_clock; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_reset; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@46401.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_io_portEnable; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  STORE_ADDR_PORT_LSQ_E_1_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@46401.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_E_1_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@46401.4]
  wire  storeEmpty; // @[LSQBRAM.scala 46:24:@46330.4 LSQBRAM.scala 151:14:@46747.4]
  wire  loadEmpty; // @[LSQBRAM.scala 52:23:@46336.4 LSQBRAM.scala 119:13:@46602.4]
  wire [1:0] bbNumStores; // @[LSQBRAM.scala 43:25:@46327.4 LSQBRAM.scala 96:15:@46487.4]
  wire [15:0] storeTail; // @[LSQBRAM.scala 44:23:@46328.4 LSQBRAM.scala 149:13:@46745.4]
  wire [15:0] storeHead; // @[LSQBRAM.scala 45:23:@46329.4 LSQBRAM.scala 150:13:@46746.4]
  wire [15:0] loadTail; // @[LSQBRAM.scala 50:22:@46334.4 LSQBRAM.scala 117:12:@46600.4]
  wire [15:0] loadHead; // @[LSQBRAM.scala 51:22:@46335.4 LSQBRAM.scala 118:12:@46601.4]
  STORE_QUEUE_LSQ_E storeQ ( // @[LSQBRAM.scala 72:22:@46354.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(storeQ_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(storeQ_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(storeQ_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(storeQ_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(storeQ_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(storeQ_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(storeQ_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(storeQ_io_bbStoreOffsets_15),
    .io_bbStorePorts_0(storeQ_io_bbStorePorts_0),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadAddressDone_8(storeQ_io_loadAddressDone_8),
    .io_loadAddressDone_9(storeQ_io_loadAddressDone_9),
    .io_loadAddressDone_10(storeQ_io_loadAddressDone_10),
    .io_loadAddressDone_11(storeQ_io_loadAddressDone_11),
    .io_loadAddressDone_12(storeQ_io_loadAddressDone_12),
    .io_loadAddressDone_13(storeQ_io_loadAddressDone_13),
    .io_loadAddressDone_14(storeQ_io_loadAddressDone_14),
    .io_loadAddressDone_15(storeQ_io_loadAddressDone_15),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadDataDone_8(storeQ_io_loadDataDone_8),
    .io_loadDataDone_9(storeQ_io_loadDataDone_9),
    .io_loadDataDone_10(storeQ_io_loadDataDone_10),
    .io_loadDataDone_11(storeQ_io_loadDataDone_11),
    .io_loadDataDone_12(storeQ_io_loadDataDone_12),
    .io_loadDataDone_13(storeQ_io_loadDataDone_13),
    .io_loadDataDone_14(storeQ_io_loadDataDone_14),
    .io_loadDataDone_15(storeQ_io_loadDataDone_15),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_loadAddressQueue_8(storeQ_io_loadAddressQueue_8),
    .io_loadAddressQueue_9(storeQ_io_loadAddressQueue_9),
    .io_loadAddressQueue_10(storeQ_io_loadAddressQueue_10),
    .io_loadAddressQueue_11(storeQ_io_loadAddressQueue_11),
    .io_loadAddressQueue_12(storeQ_io_loadAddressQueue_12),
    .io_loadAddressQueue_13(storeQ_io_loadAddressQueue_13),
    .io_loadAddressQueue_14(storeQ_io_loadAddressQueue_14),
    .io_loadAddressQueue_15(storeQ_io_loadAddressQueue_15),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(storeQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(storeQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(storeQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(storeQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(storeQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(storeQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(storeQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(storeQ_io_storeAddrDone_15),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeDataDone_8(storeQ_io_storeDataDone_8),
    .io_storeDataDone_9(storeQ_io_storeDataDone_9),
    .io_storeDataDone_10(storeQ_io_storeDataDone_10),
    .io_storeDataDone_11(storeQ_io_storeDataDone_11),
    .io_storeDataDone_12(storeQ_io_storeDataDone_12),
    .io_storeDataDone_13(storeQ_io_storeDataDone_13),
    .io_storeDataDone_14(storeQ_io_storeDataDone_14),
    .io_storeDataDone_15(storeQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(storeQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(storeQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(storeQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(storeQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(storeQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(storeQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(storeQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(storeQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(storeQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(storeQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(storeQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(storeQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(storeQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(storeQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(storeQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(storeQ_io_storeDataQueue_15),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_storeDataEnable_1(storeQ_io_storeDataEnable_1),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_dataFromStorePorts_1(storeQ_io_dataFromStorePorts_1),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_storeAddrEnable_1(storeQ_io_storeAddrEnable_1),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_addressFromStorePorts_1(storeQ_io_addressFromStorePorts_1),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeEnableToMem(storeQ_io_storeEnableToMem),
    .io_memIsReadyForStores(storeQ_io_memIsReadyForStores)
  );
  LOAD_QUEUE_LSQ_E loadQ ( // @[LSQBRAM.scala 73:21:@46357.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(loadQ_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(loadQ_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(loadQ_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(loadQ_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(loadQ_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(loadQ_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(loadQ_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(loadQ_io_bbLoadOffsets_15),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(loadQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(loadQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(loadQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(loadQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(loadQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(loadQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(loadQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(loadQ_io_storeAddrDone_15),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeDataDone_8(loadQ_io_storeDataDone_8),
    .io_storeDataDone_9(loadQ_io_storeDataDone_9),
    .io_storeDataDone_10(loadQ_io_storeDataDone_10),
    .io_storeDataDone_11(loadQ_io_storeDataDone_11),
    .io_storeDataDone_12(loadQ_io_storeDataDone_12),
    .io_storeDataDone_13(loadQ_io_storeDataDone_13),
    .io_storeDataDone_14(loadQ_io_storeDataDone_14),
    .io_storeDataDone_15(loadQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(loadQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(loadQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(loadQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(loadQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(loadQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(loadQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(loadQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(loadQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(loadQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(loadQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(loadQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(loadQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(loadQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(loadQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(loadQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(loadQ_io_storeDataQueue_15),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadAddrDone_8(loadQ_io_loadAddrDone_8),
    .io_loadAddrDone_9(loadQ_io_loadAddrDone_9),
    .io_loadAddrDone_10(loadQ_io_loadAddrDone_10),
    .io_loadAddrDone_11(loadQ_io_loadAddrDone_11),
    .io_loadAddrDone_12(loadQ_io_loadAddrDone_12),
    .io_loadAddrDone_13(loadQ_io_loadAddrDone_13),
    .io_loadAddrDone_14(loadQ_io_loadAddrDone_14),
    .io_loadAddrDone_15(loadQ_io_loadAddrDone_15),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadDataDone_8(loadQ_io_loadDataDone_8),
    .io_loadDataDone_9(loadQ_io_loadDataDone_9),
    .io_loadDataDone_10(loadQ_io_loadDataDone_10),
    .io_loadDataDone_11(loadQ_io_loadDataDone_11),
    .io_loadDataDone_12(loadQ_io_loadDataDone_12),
    .io_loadDataDone_13(loadQ_io_loadDataDone_13),
    .io_loadDataDone_14(loadQ_io_loadDataDone_14),
    .io_loadDataDone_15(loadQ_io_loadDataDone_15),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrQueue_8(loadQ_io_loadAddrQueue_8),
    .io_loadAddrQueue_9(loadQ_io_loadAddrQueue_9),
    .io_loadAddrQueue_10(loadQ_io_loadAddrQueue_10),
    .io_loadAddrQueue_11(loadQ_io_loadAddrQueue_11),
    .io_loadAddrQueue_12(loadQ_io_loadAddrQueue_12),
    .io_loadAddrQueue_13(loadQ_io_loadAddrQueue_13),
    .io_loadAddrQueue_14(loadQ_io_loadAddrQueue_14),
    .io_loadAddrQueue_15(loadQ_io_loadAddrQueue_15),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadEnableToMem(loadQ_io_loadEnableToMem),
    .io_memIsReadyForLoads(loadQ_io_memIsReadyForLoads)
  );
  GROUP_ALLOCATOR_LSQ_E GA ( // @[LSQBRAM.scala 74:18:@46360.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(GA_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(GA_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(GA_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(GA_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(GA_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(GA_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(GA_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(GA_io_bbLoadOffsets_15),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(GA_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(GA_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(GA_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(GA_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(GA_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(GA_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(GA_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(GA_io_bbStoreOffsets_15),
    .io_bbStorePorts_0(GA_io_bbStorePorts_0),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_bbStartSignals_1(GA_io_bbStartSignals_1),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_readyToPrevious_1(GA_io_readyToPrevious_1),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0),
    .io_storePortsEnable_1(GA_io_storePortsEnable_1)
  );
  LOAD_PORT_LSQ_E LOAD_PORT_LSQ_E ( // @[LSQBRAM.scala 77:11:@46363.4]
    .clock(LOAD_PORT_LSQ_E_clock),
    .reset(LOAD_PORT_LSQ_E_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_E_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_E_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_E_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_E_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_E_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_E_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_E_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_E_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_E_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_E_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_E_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_E_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_E STORE_DATA_PORT_LSQ_E ( // @[LSQBRAM.scala 80:11:@46379.4]
    .clock(STORE_DATA_PORT_LSQ_E_clock),
    .reset(STORE_DATA_PORT_LSQ_E_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_E_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_E_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_E_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_E_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_E_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_E_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_E STORE_DATA_PORT_LSQ_E_1 ( // @[LSQBRAM.scala 80:11:@46382.4]
    .clock(STORE_DATA_PORT_LSQ_E_1_clock),
    .reset(STORE_DATA_PORT_LSQ_E_1_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_E_1_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_E_1_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_E_1_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_E STORE_ADDR_PORT_LSQ_E ( // @[LSQBRAM.scala 83:11:@46398.4]
    .clock(STORE_ADDR_PORT_LSQ_E_clock),
    .reset(STORE_ADDR_PORT_LSQ_E_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_E_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_E_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_E_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_E STORE_ADDR_PORT_LSQ_E_1 ( // @[LSQBRAM.scala 83:11:@46401.4]
    .clock(STORE_ADDR_PORT_LSQ_E_1_clock),
    .reset(STORE_ADDR_PORT_LSQ_E_1_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_E_1_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_E_1_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_E_1_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 46:24:@46330.4 LSQBRAM.scala 151:14:@46747.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 52:23:@46336.4 LSQBRAM.scala 119:13:@46602.4]
  assign bbNumStores = GA_io_bbNumStores; // @[LSQBRAM.scala 43:25:@46327.4 LSQBRAM.scala 96:15:@46487.4]
  assign storeTail = {{12'd0}, storeQ_io_storeTail}; // @[LSQBRAM.scala 44:23:@46328.4 LSQBRAM.scala 149:13:@46745.4]
  assign storeHead = {{12'd0}, storeQ_io_storeHead}; // @[LSQBRAM.scala 45:23:@46329.4 LSQBRAM.scala 150:13:@46746.4]
  assign loadTail = {{12'd0}, loadQ_io_loadTail}; // @[LSQBRAM.scala 50:22:@46334.4 LSQBRAM.scala 117:12:@46600.4]
  assign loadHead = {{12'd0}, loadQ_io_loadHead}; // @[LSQBRAM.scala 51:22:@46335.4 LSQBRAM.scala 118:12:@46601.4]
  assign io_storeDataOut = storeQ_io_storeDataToMem; // @[LSQBRAM.scala 161:19:@46821.4]
  assign io_storeAddrOut = storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 160:19:@46820.4]
  assign io_storeEnable = storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 162:18:@46822.4]
  assign io_loadAddrOut = loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 135:18:@46658.4]
  assign io_loadEnable = loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 136:17:@46659.4]
  assign io_bbReadyToPrevs_0 = GA_io_readyToPrevious_0; // @[LSQBRAM.scala 102:21:@46494.4]
  assign io_bbReadyToPrevs_1 = GA_io_readyToPrevious_1; // @[LSQBRAM.scala 102:21:@46495.4]
  assign io_rdPortsPrev_0_ready = LOAD_PORT_LSQ_E_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@46826.4]
  assign io_rdPortsNext_0_valid = LOAD_PORT_LSQ_E_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@46829.4]
  assign io_rdPortsNext_0_bits = LOAD_PORT_LSQ_E_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@46828.4]
  assign io_wrAddrPorts_0_ready = STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@46844.4]
  assign io_wrAddrPorts_1_ready = STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@46856.4]
  assign io_wrDataPorts_0_ready = STORE_DATA_PORT_LSQ_E_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@46838.4]
  assign io_wrDataPorts_1_ready = STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@46850.4]
  assign io_Empty_Valid = storeEmpty & loadEmpty; // @[LSQBRAM.scala 86:18:@46418.4]
  assign storeQ_clock = clock; // @[:@46355.4]
  assign storeQ_reset = reset; // @[:@46356.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 145:21:@46711.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 146:28:@46712.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 146:28:@46713.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 146:28:@46714.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 146:28:@46715.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 146:28:@46716.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 146:28:@46717.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 146:28:@46718.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 146:28:@46719.4]
  assign storeQ_io_bbStoreOffsets_8 = GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 146:28:@46720.4]
  assign storeQ_io_bbStoreOffsets_9 = GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 146:28:@46721.4]
  assign storeQ_io_bbStoreOffsets_10 = GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 146:28:@46722.4]
  assign storeQ_io_bbStoreOffsets_11 = GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 146:28:@46723.4]
  assign storeQ_io_bbStoreOffsets_12 = GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 146:28:@46724.4]
  assign storeQ_io_bbStoreOffsets_13 = GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 146:28:@46725.4]
  assign storeQ_io_bbStoreOffsets_14 = GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 146:28:@46726.4]
  assign storeQ_io_bbStoreOffsets_15 = GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 146:28:@46727.4]
  assign storeQ_io_bbStorePorts_0 = GA_io_bbStorePorts_0; // @[LSQBRAM.scala 147:26:@46728.4]
  assign storeQ_io_bbNumStores = bbNumStores[0]; // @[LSQBRAM.scala 148:25:@46744.4]
  assign storeQ_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 139:22:@46660.4]
  assign storeQ_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 140:22:@46661.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 141:23:@46662.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 142:29:@46663.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 142:29:@46664.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 142:29:@46665.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 142:29:@46666.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 142:29:@46667.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 142:29:@46668.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 142:29:@46669.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 142:29:@46670.4]
  assign storeQ_io_loadAddressDone_8 = loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 142:29:@46671.4]
  assign storeQ_io_loadAddressDone_9 = loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 142:29:@46672.4]
  assign storeQ_io_loadAddressDone_10 = loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 142:29:@46673.4]
  assign storeQ_io_loadAddressDone_11 = loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 142:29:@46674.4]
  assign storeQ_io_loadAddressDone_12 = loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 142:29:@46675.4]
  assign storeQ_io_loadAddressDone_13 = loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 142:29:@46676.4]
  assign storeQ_io_loadAddressDone_14 = loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 142:29:@46677.4]
  assign storeQ_io_loadAddressDone_15 = loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 142:29:@46678.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 143:26:@46679.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 143:26:@46680.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 143:26:@46681.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 143:26:@46682.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 143:26:@46683.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 143:26:@46684.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 143:26:@46685.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 143:26:@46686.4]
  assign storeQ_io_loadDataDone_8 = loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 143:26:@46687.4]
  assign storeQ_io_loadDataDone_9 = loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 143:26:@46688.4]
  assign storeQ_io_loadDataDone_10 = loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 143:26:@46689.4]
  assign storeQ_io_loadDataDone_11 = loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 143:26:@46690.4]
  assign storeQ_io_loadDataDone_12 = loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 143:26:@46691.4]
  assign storeQ_io_loadDataDone_13 = loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 143:26:@46692.4]
  assign storeQ_io_loadDataDone_14 = loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 143:26:@46693.4]
  assign storeQ_io_loadDataDone_15 = loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 143:26:@46694.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 144:30:@46695.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 144:30:@46696.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 144:30:@46697.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 144:30:@46698.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 144:30:@46699.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 144:30:@46700.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 144:30:@46701.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 144:30:@46702.4]
  assign storeQ_io_loadAddressQueue_8 = loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 144:30:@46703.4]
  assign storeQ_io_loadAddressQueue_9 = loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 144:30:@46704.4]
  assign storeQ_io_loadAddressQueue_10 = loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 144:30:@46705.4]
  assign storeQ_io_loadAddressQueue_11 = loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 144:30:@46706.4]
  assign storeQ_io_loadAddressQueue_12 = loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 144:30:@46707.4]
  assign storeQ_io_loadAddressQueue_13 = loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 144:30:@46708.4]
  assign storeQ_io_loadAddressQueue_14 = loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 144:30:@46709.4]
  assign storeQ_io_loadAddressQueue_15 = loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 144:30:@46710.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_E_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@46812.4]
  assign storeQ_io_storeDataEnable_1 = STORE_DATA_PORT_LSQ_E_1_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@46813.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_E_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@46814.4]
  assign storeQ_io_dataFromStorePorts_1 = STORE_DATA_PORT_LSQ_E_1_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@46815.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_E_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@46816.4]
  assign storeQ_io_storeAddrEnable_1 = STORE_ADDR_PORT_LSQ_E_1_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@46817.4]
  assign storeQ_io_addressFromStorePorts_0 = STORE_ADDR_PORT_LSQ_E_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@46818.4]
  assign storeQ_io_addressFromStorePorts_1 = STORE_ADDR_PORT_LSQ_E_1_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@46819.4]
  assign storeQ_io_memIsReadyForStores = io_memIsReadyForStores; // @[LSQBRAM.scala 163:33:@46823.4]
  assign loadQ_clock = clock; // @[:@46358.4]
  assign loadQ_reset = reset; // @[:@46359.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 113:20:@46566.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 114:26:@46567.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 114:26:@46568.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 114:26:@46569.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 114:26:@46570.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 114:26:@46571.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 114:26:@46572.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 114:26:@46573.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 114:26:@46574.4]
  assign loadQ_io_bbLoadOffsets_8 = GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 114:26:@46575.4]
  assign loadQ_io_bbLoadOffsets_9 = GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 114:26:@46576.4]
  assign loadQ_io_bbLoadOffsets_10 = GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 114:26:@46577.4]
  assign loadQ_io_bbLoadOffsets_11 = GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 114:26:@46578.4]
  assign loadQ_io_bbLoadOffsets_12 = GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 114:26:@46579.4]
  assign loadQ_io_bbLoadOffsets_13 = GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 114:26:@46580.4]
  assign loadQ_io_bbLoadOffsets_14 = GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 114:26:@46581.4]
  assign loadQ_io_bbLoadOffsets_15 = GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 114:26:@46582.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQBRAM.scala 116:23:@46599.4]
  assign loadQ_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 106:22:@46499.4]
  assign loadQ_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 107:22:@46500.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 108:23:@46501.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 109:26:@46502.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 109:26:@46503.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 109:26:@46504.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 109:26:@46505.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 109:26:@46506.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 109:26:@46507.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 109:26:@46508.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 109:26:@46509.4]
  assign loadQ_io_storeAddrDone_8 = storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 109:26:@46510.4]
  assign loadQ_io_storeAddrDone_9 = storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 109:26:@46511.4]
  assign loadQ_io_storeAddrDone_10 = storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 109:26:@46512.4]
  assign loadQ_io_storeAddrDone_11 = storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 109:26:@46513.4]
  assign loadQ_io_storeAddrDone_12 = storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 109:26:@46514.4]
  assign loadQ_io_storeAddrDone_13 = storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 109:26:@46515.4]
  assign loadQ_io_storeAddrDone_14 = storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 109:26:@46516.4]
  assign loadQ_io_storeAddrDone_15 = storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 109:26:@46517.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 110:26:@46518.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 110:26:@46519.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 110:26:@46520.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 110:26:@46521.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 110:26:@46522.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 110:26:@46523.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 110:26:@46524.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 110:26:@46525.4]
  assign loadQ_io_storeDataDone_8 = storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 110:26:@46526.4]
  assign loadQ_io_storeDataDone_9 = storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 110:26:@46527.4]
  assign loadQ_io_storeDataDone_10 = storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 110:26:@46528.4]
  assign loadQ_io_storeDataDone_11 = storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 110:26:@46529.4]
  assign loadQ_io_storeDataDone_12 = storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 110:26:@46530.4]
  assign loadQ_io_storeDataDone_13 = storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 110:26:@46531.4]
  assign loadQ_io_storeDataDone_14 = storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 110:26:@46532.4]
  assign loadQ_io_storeDataDone_15 = storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 110:26:@46533.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 111:27:@46534.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 111:27:@46535.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 111:27:@46536.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 111:27:@46537.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 111:27:@46538.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 111:27:@46539.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 111:27:@46540.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 111:27:@46541.4]
  assign loadQ_io_storeAddrQueue_8 = storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 111:27:@46542.4]
  assign loadQ_io_storeAddrQueue_9 = storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 111:27:@46543.4]
  assign loadQ_io_storeAddrQueue_10 = storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 111:27:@46544.4]
  assign loadQ_io_storeAddrQueue_11 = storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 111:27:@46545.4]
  assign loadQ_io_storeAddrQueue_12 = storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 111:27:@46546.4]
  assign loadQ_io_storeAddrQueue_13 = storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 111:27:@46547.4]
  assign loadQ_io_storeAddrQueue_14 = storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 111:27:@46548.4]
  assign loadQ_io_storeAddrQueue_15 = storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 111:27:@46549.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 112:27:@46550.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 112:27:@46551.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 112:27:@46552.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 112:27:@46553.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 112:27:@46554.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 112:27:@46555.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 112:27:@46556.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 112:27:@46557.4]
  assign loadQ_io_storeDataQueue_8 = storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 112:27:@46558.4]
  assign loadQ_io_storeDataQueue_9 = storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 112:27:@46559.4]
  assign loadQ_io_storeDataQueue_10 = storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 112:27:@46560.4]
  assign loadQ_io_storeDataQueue_11 = storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 112:27:@46561.4]
  assign loadQ_io_storeDataQueue_12 = storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 112:27:@46562.4]
  assign loadQ_io_storeDataQueue_13 = storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 112:27:@46563.4]
  assign loadQ_io_storeDataQueue_14 = storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 112:27:@46564.4]
  assign loadQ_io_storeDataQueue_15 = storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 112:27:@46565.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_E_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@46655.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_E_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@46654.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_E_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@46653.4]
  assign loadQ_io_loadDataFromMem = io_loadDataIn; // @[LSQBRAM.scala 133:28:@46656.4]
  assign loadQ_io_memIsReadyForLoads = io_memIsReadyForLoads; // @[LSQBRAM.scala 134:31:@46657.4]
  assign GA_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 91:18:@46452.4]
  assign GA_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 92:18:@46453.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 93:19:@46454.4]
  assign GA_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 97:19:@46488.4]
  assign GA_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 98:19:@46489.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 99:20:@46490.4]
  assign GA_io_bbStartSignals_0 = io_bbpValids_0; // @[LSQBRAM.scala 101:24:@46492.4]
  assign GA_io_bbStartSignals_1 = io_bbpValids_1; // @[LSQBRAM.scala 101:24:@46493.4]
  assign LOAD_PORT_LSQ_E_clock = clock; // @[:@46364.4]
  assign LOAD_PORT_LSQ_E_reset = reset; // @[:@46365.4]
  assign LOAD_PORT_LSQ_E_io_addrFromPrev_valid = io_rdPortsPrev_0_valid; // @[LSQBRAM.scala 76:26:@46377.4]
  assign LOAD_PORT_LSQ_E_io_addrFromPrev_bits = io_rdPortsPrev_0_bits; // @[LSQBRAM.scala 76:26:@46376.4]
  assign LOAD_PORT_LSQ_E_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 76:26:@46375.4]
  assign LOAD_PORT_LSQ_E_io_dataToNext_ready = io_rdPortsNext_0_ready; // @[LSQBRAM.scala 76:26:@46374.4]
  assign LOAD_PORT_LSQ_E_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 76:26:@46368.4]
  assign LOAD_PORT_LSQ_E_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 76:26:@46367.4]
  assign STORE_DATA_PORT_LSQ_E_clock = clock; // @[:@46380.4]
  assign STORE_DATA_PORT_LSQ_E_reset = reset; // @[:@46381.4]
  assign STORE_DATA_PORT_LSQ_E_io_dataFromPrev_valid = io_wrDataPorts_0_valid; // @[LSQBRAM.scala 79:31:@46390.4]
  assign STORE_DATA_PORT_LSQ_E_io_dataFromPrev_bits = io_wrDataPorts_0_bits; // @[LSQBRAM.scala 79:31:@46389.4]
  assign STORE_DATA_PORT_LSQ_E_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 79:31:@46388.4]
  assign STORE_DATA_PORT_LSQ_E_1_clock = clock; // @[:@46383.4]
  assign STORE_DATA_PORT_LSQ_E_1_reset = reset; // @[:@46384.4]
  assign STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_valid = io_wrDataPorts_1_valid; // @[LSQBRAM.scala 79:31:@46396.4]
  assign STORE_DATA_PORT_LSQ_E_1_io_dataFromPrev_bits = io_wrDataPorts_1_bits; // @[LSQBRAM.scala 79:31:@46395.4]
  assign STORE_DATA_PORT_LSQ_E_1_io_portEnable = GA_io_storePortsEnable_1; // @[LSQBRAM.scala 79:31:@46394.4]
  assign STORE_ADDR_PORT_LSQ_E_clock = clock; // @[:@46399.4]
  assign STORE_ADDR_PORT_LSQ_E_reset = reset; // @[:@46400.4]
  assign STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_valid = io_wrAddrPorts_0_valid; // @[LSQBRAM.scala 82:34:@46409.4]
  assign STORE_ADDR_PORT_LSQ_E_io_dataFromPrev_bits = io_wrAddrPorts_0_bits; // @[LSQBRAM.scala 82:34:@46408.4]
  assign STORE_ADDR_PORT_LSQ_E_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 82:34:@46407.4]
  assign STORE_ADDR_PORT_LSQ_E_1_clock = clock; // @[:@46402.4]
  assign STORE_ADDR_PORT_LSQ_E_1_reset = reset; // @[:@46403.4]
  assign STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_valid = io_wrAddrPorts_1_valid; // @[LSQBRAM.scala 82:34:@46415.4]
  assign STORE_ADDR_PORT_LSQ_E_1_io_dataFromPrev_bits = io_wrAddrPorts_1_bits; // @[LSQBRAM.scala 82:34:@46414.4]
  assign STORE_ADDR_PORT_LSQ_E_1_io_portEnable = GA_io_storePortsEnable_1; // @[LSQBRAM.scala 82:34:@46413.4]
endmodule
