// tb.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module tb (
	);

	wire  [255:0] if_loop_3_inst_avmm_1_rw_readdata;                                                           // mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_readdata -> if_loop_3_inst:avmm_1_rw_readdata
	wire   [31:0] if_loop_3_inst_avmm_1_rw_address;                                                            // if_loop_3_inst:avmm_1_rw_address -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_address
	wire   [31:0] if_loop_3_inst_avmm_1_rw_byteenable;                                                         // if_loop_3_inst:avmm_1_rw_byteenable -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_byteenable
	wire          if_loop_3_inst_avmm_1_rw_read;                                                               // if_loop_3_inst:avmm_1_rw_read -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_read
	wire          if_loop_3_inst_avmm_1_rw_write;                                                              // if_loop_3_inst:avmm_1_rw_write -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_write
	wire  [255:0] if_loop_3_inst_avmm_1_rw_writedata;                                                          // if_loop_3_inst:avmm_1_rw_writedata -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:avs_writedata
	wire  [255:0] if_loop_3_inst_avmm_4_rw_readdata;                                                           // mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_readdata -> if_loop_3_inst:avmm_4_rw_readdata
	wire   [31:0] if_loop_3_inst_avmm_4_rw_address;                                                            // if_loop_3_inst:avmm_4_rw_address -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_address
	wire   [31:0] if_loop_3_inst_avmm_4_rw_byteenable;                                                         // if_loop_3_inst:avmm_4_rw_byteenable -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_byteenable
	wire          if_loop_3_inst_avmm_4_rw_read;                                                               // if_loop_3_inst:avmm_4_rw_read -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_read
	wire          if_loop_3_inst_avmm_4_rw_write;                                                              // if_loop_3_inst:avmm_4_rw_write -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_write
	wire  [255:0] if_loop_3_inst_avmm_4_rw_writedata;                                                          // if_loop_3_inst:avmm_4_rw_writedata -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:avs_writedata
	wire          clock_reset_inst_clock_clk;                                                                  // clock_reset_inst:clock -> [component_dpi_controller_if_loop_3_inst:clock, if_loop_3_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:clock, mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:clock, stream_source_dpi_bfm_if_loop_3_a_inst:clock, stream_source_dpi_bfm_if_loop_3_b_inst:clock, stream_source_dpi_bfm_if_loop_3_n_inst:clock]
	wire          clock_reset_inst_clock2x_clk;                                                                // clock_reset_inst:clock2x -> [component_dpi_controller_if_loop_3_inst:clock2x, main_dpi_controller_inst:clock2x, stream_source_dpi_bfm_if_loop_3_a_inst:clock2x, stream_source_dpi_bfm_if_loop_3_b_inst:clock2x, stream_source_dpi_bfm_if_loop_3_n_inst:clock2x]
	wire          component_dpi_controller_if_loop_3_inst_component_call_valid;                                // component_dpi_controller_if_loop_3_inst:start -> if_loop_3_inst:start
	wire          if_loop_3_inst_call_stall;                                                                   // if_loop_3_inst:busy -> component_dpi_controller_if_loop_3_inst:busy
	wire          component_dpi_controller_if_loop_3_inst_component_done_conduit;                              // component_dpi_controller_if_loop_3_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire    [0:0] main_dpi_controller_inst_component_enabled_conduit;                                          // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire          component_dpi_controller_if_loop_3_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_if_loop_3_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire          component_dpi_controller_if_loop_3_inst_dpi_control_bind_conduit;                            // component_dpi_controller_if_loop_3_inst:bind_interfaces -> if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire          component_dpi_controller_if_loop_3_inst_dpi_control_enable_conduit;                          // component_dpi_controller_if_loop_3_inst:enable_interfaces -> if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire          concatenate_component_done_inst_out_conduit_conduit;                                         // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire          concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                       // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire          split_component_start_inst_out_conduit_0_conduit;                                            // split_component_start_inst:out_conduit_0 -> component_dpi_controller_if_loop_3_inst:component_enabled
	wire          if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_if_loop_3_a_inst:do_bind
	wire          if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_if_loop_3_a_inst:enable
	wire          if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_if_loop_3_a_inst:source_ready
	wire          if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:do_bind
	wire          if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:enable
	wire          if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> stream_source_dpi_bfm_if_loop_3_b_inst:source_ready
	wire          if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit;           // if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_2 -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:do_bind
	wire          if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit;         // if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_2 -> mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:enable
	wire          if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit; // if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_2 -> stream_source_dpi_bfm_if_loop_3_n_inst:source_ready
	wire          if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit;           // if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_if_loop_3_b_inst:do_bind
	wire          if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit;         // if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_3 -> stream_source_dpi_bfm_if_loop_3_b_inst:enable
	wire          if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit;           // if_loop_3_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_if_loop_3_n_inst:do_bind
	wire          if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit;         // if_loop_3_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_4 -> stream_source_dpi_bfm_if_loop_3_n_inst:enable
	wire          component_dpi_controller_if_loop_3_inst_read_implicit_streams_conduit;                       // component_dpi_controller_if_loop_3_inst:read_implicit_streams -> if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire          main_dpi_controller_inst_reset_ctrl_conduit;                                                 // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire          if_loop_3_inst_return_valid;                                                                 // if_loop_3_inst:done -> component_dpi_controller_if_loop_3_inst:done
	wire          component_dpi_controller_if_loop_3_inst_component_return_stall;                              // component_dpi_controller_if_loop_3_inst:stall -> if_loop_3_inst:stall
	wire   [31:0] if_loop_3_inst_returndata_data;                                                              // if_loop_3_inst:returndata -> component_dpi_controller_if_loop_3_inst:returndata
	wire   [63:0] stream_source_dpi_bfm_if_loop_3_a_inst_source_data_data;                                     // stream_source_dpi_bfm_if_loop_3_a_inst:source_data -> if_loop_3_inst:a
	wire   [63:0] stream_source_dpi_bfm_if_loop_3_b_inst_source_data_data;                                     // stream_source_dpi_bfm_if_loop_3_b_inst:source_data -> if_loop_3_inst:b
	wire   [31:0] stream_source_dpi_bfm_if_loop_3_n_inst_source_data_data;                                     // stream_source_dpi_bfm_if_loop_3_n_inst:source_data -> if_loop_3_inst:n
	wire          clock_reset_inst_reset_reset;                                                                // clock_reset_inst:resetn -> [component_dpi_controller_if_loop_3_inst:resetn, if_loop_3_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst:reset_n, mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst:reset_n, stream_source_dpi_bfm_if_loop_3_a_inst:resetn, stream_source_dpi_bfm_if_loop_3_b_inst:resetn, stream_source_dpi_bfm_if_loop_3_n_inst:resetn]
	wire          component_dpi_controller_if_loop_3_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_if_loop_3_inst:done_irq

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("if_loop_3"),
		.COMPONENT_MANGLED_NAME       ("\\3fif_loop_3@@YAHAEAV\\3f$mm_host@HU\\3f$dwidth@$0BAA@@ihc@@U\\3f$awidth@$0CA@@2@U\\3f$aspace@$00@2@U\\3f$latency@$00@2@@ihc@@AEAV\\3f$mm_host@HU\\3f$dwidth@$0BAA@@ihc@@U\\3f$awidth@$0CA@@2@U\\3f$aspace@$03@2@U\\3f$latency@$00@2@@2@H@Z"),
		.RETURN_DATAWIDTH             (32),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_if_loop_3_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                       //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                     //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                     //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_if_loop_3_inst_dpi_control_bind_conduit),                 //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_if_loop_3_inst_dpi_control_enable_conduit),               //               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                 //                component_enabled.conduit
		.component_done                   (component_dpi_controller_if_loop_3_inst_component_done_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_if_loop_3_inst_component_wait_for_stream_writes_conduit), // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                                 //                       agent_busy.conduit
		.read_implicit_streams            (component_dpi_controller_if_loop_3_inst_read_implicit_streams_conduit),            //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                                 //             readback_from_agents.conduit
		.start                            (component_dpi_controller_if_loop_3_inst_component_call_valid),                     //                   component_call.valid
		.busy                             (if_loop_3_inst_call_stall),                                                        //                                 .stall
		.done                             (if_loop_3_inst_return_valid),                                                      //                 component_return.valid
		.stall                            (component_dpi_controller_if_loop_3_inst_component_return_stall),                   //                                 .stall
		.done_irq                         (component_dpi_controller_if_loop_3_inst_component_irq_irq),                        //                    component_irq.irq
		.returndata                       (if_loop_3_inst_returndata_data)                                                    //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),            //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_if_loop_3_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),            //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_if_loop_3_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	tb_if_loop_3_component_dpi_controller_bind_conduit_fanout_inst if_loop_3_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_if_loop_3_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_if_loop_3_component_dpi_controller_bind_conduit_fanout_inst if_loop_3_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_if_loop_3_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // out_conduit_2.conduit
		.out_conduit_3 (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit), // out_conduit_3.conduit
		.out_conduit_4 (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit)  // out_conduit_4.conduit
	);

	tb_if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_if_loop_3_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), // out_conduit_1.conduit
		.out_conduit_2 (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit)  // out_conduit_2.conduit
	);

	tb_if_loop_3_inst if_loop_3_inst (
		.a                    (stream_source_dpi_bfm_if_loop_3_a_inst_source_data_data),        //          a.data
		.avmm_1_rw_address    (if_loop_3_inst_avmm_1_rw_address),                               //  avmm_1_rw.address
		.avmm_1_rw_byteenable (if_loop_3_inst_avmm_1_rw_byteenable),                            //           .byteenable
		.avmm_1_rw_read       (if_loop_3_inst_avmm_1_rw_read),                                  //           .read
		.avmm_1_rw_readdata   (if_loop_3_inst_avmm_1_rw_readdata),                              //           .readdata
		.avmm_1_rw_write      (if_loop_3_inst_avmm_1_rw_write),                                 //           .write
		.avmm_1_rw_writedata  (if_loop_3_inst_avmm_1_rw_writedata),                             //           .writedata
		.avmm_4_rw_address    (if_loop_3_inst_avmm_4_rw_address),                               //  avmm_4_rw.address
		.avmm_4_rw_byteenable (if_loop_3_inst_avmm_4_rw_byteenable),                            //           .byteenable
		.avmm_4_rw_read       (if_loop_3_inst_avmm_4_rw_read),                                  //           .read
		.avmm_4_rw_readdata   (if_loop_3_inst_avmm_4_rw_readdata),                              //           .readdata
		.avmm_4_rw_write      (if_loop_3_inst_avmm_4_rw_write),                                 //           .write
		.avmm_4_rw_writedata  (if_loop_3_inst_avmm_4_rw_writedata),                             //           .writedata
		.b                    (stream_source_dpi_bfm_if_loop_3_b_inst_source_data_data),        //          b.data
		.start                (component_dpi_controller_if_loop_3_inst_component_call_valid),   //       call.valid
		.busy                 (if_loop_3_inst_call_stall),                                      //           .stall
		.clock                (clock_reset_inst_clock_clk),                                     //      clock.clk
		.n                    (stream_source_dpi_bfm_if_loop_3_n_inst_source_data_data),        //          n.data
		.resetn               (clock_reset_inst_reset_reset),                                   //      reset.reset_n
		.done                 (if_loop_3_inst_return_valid),                                    //     return.valid
		.stall                (component_dpi_controller_if_loop_3_inst_component_return_stall), //           .stall
		.returndata           (if_loop_3_inst_returndata_data)                                  // returndata.data
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (1),
		.COMPONENT_NAMES_STR ("if_loop_3")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (32),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("if_loop_3"),
		.INTERFACE_ID               (1)
	) mm_agent_dpi_bfm_if_loop_3_avmm_1_rw_inst (
		.do_bind           (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),   //   dpi_control_bind.conduit
		.enable            (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                          //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                        //              reset.reset_n
		.avs_writedata     (if_loop_3_inst_avmm_1_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (if_loop_3_inst_avmm_1_rw_readdata),                                                   //                   .readdata
		.avs_address       (if_loop_3_inst_avmm_1_rw_address),                                                    //                   .address
		.avs_write         (if_loop_3_inst_avmm_1_rw_write),                                                      //                   .write
		.avs_read          (if_loop_3_inst_avmm_1_rw_read),                                                       //                   .read
		.avs_byteenable    (if_loop_3_inst_avmm_1_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                     //        (terminated)
	);

	hls_sim_mm_agent_dpi_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (32),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.COMPONENT_NAME             ("if_loop_3"),
		.INTERFACE_ID               (4)
	) mm_agent_dpi_bfm_if_loop_3_avmm_4_rw_inst (
		.do_bind           (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_2_conduit),   //   dpi_control_bind.conduit
		.enable            (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_2_conduit), // dpi_control_enable.conduit
		.clock             (clock_reset_inst_clock_clk),                                                          //              clock.clk
		.reset_n           (clock_reset_inst_reset_reset),                                                        //              reset.reset_n
		.avs_writedata     (if_loop_3_inst_avmm_4_rw_writedata),                                                  //                 s0.writedata
		.avs_readdata      (if_loop_3_inst_avmm_4_rw_readdata),                                                   //                   .readdata
		.avs_address       (if_loop_3_inst_avmm_4_rw_address),                                                    //                   .address
		.avs_write         (if_loop_3_inst_avmm_4_rw_write),                                                      //                   .write
		.avs_read          (if_loop_3_inst_avmm_4_rw_read),                                                       //                   .read
		.avs_byteenable    (if_loop_3_inst_avmm_4_rw_byteenable),                                                 //                   .byteenable
		.avs_readdatavalid ()                                                                                     //        (terminated)
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("if_loop_3"),
		.INTERFACE_NAME                  ("a"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_if_loop_3_a_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                  //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                //            clock2x.clk
		.do_bind      (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //   dpi_control_bind.conduit
		.enable       (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_if_loop_3_a_inst_source_data_data),                                     //        source_data.data
		.source_ready (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //       source_ready.conduit
		.source_valid ()                                                                                             //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("if_loop_3"),
		.INTERFACE_NAME                  ("b"),
		.STREAM_DATAWIDTH                (64),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_if_loop_3_b_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                  //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                //            clock2x.clk
		.do_bind      (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_3_conduit),           //   dpi_control_bind.conduit
		.enable       (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_3_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_if_loop_3_b_inst_source_data_data),                                     //        source_data.data
		.source_ready (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //       source_ready.conduit
		.source_valid ()                                                                                             //             source.conduit
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("if_loop_3"),
		.INTERFACE_NAME                  ("n"),
		.STREAM_DATAWIDTH                (32),
		.STREAM_BITSPERSYMBOL            (1),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_if_loop_3_n_inst (
		.clock        (clock_reset_inst_clock_clk),                                                                  //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                                //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                                //            clock2x.clk
		.do_bind      (if_loop_3_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_4_conduit),           //   dpi_control_bind.conduit
		.enable       (if_loop_3_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_4_conduit),         // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_if_loop_3_n_inst_source_data_data),                                     //        source_data.data
		.source_ready (if_loop_3_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_2_conduit), //       source_ready.conduit
		.source_valid ()                                                                                             //             source.conduit
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                                //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                             // clk_reset.reset
		.sender_irq (component_dpi_controller_if_loop_3_inst_component_irq_irq)  //    sender.irq
	);

endmodule
