`ifndef _DDR5MC_BFM_NA_NOC_REGS_DEFINES_VH_
`define _DDR5MC_BFM_NA_NOC_REGS_DEFINES_VH_

// spyglass disable_block ConstName
/* Address and Field defines*/

/* PCSR_LOCK */
`define DDRMC5_NOC_PCSR_LOCK_OFFSET 17'hc
`define DDRMC5_NOC_PCSR_LOCK_FLD_STATE 0
`define DDRMC5_NOC_PCSR_LOCK_FLD_STATE_WIDTH 1
`define DDRMC5_NOC_PCSR_LOCK_FLD_RESERVED 31:1
`define DDRMC5_NOC_PCSR_LOCK_FLD_RESERVED_WIDTH 31
`define DDRMC5_NOC_PCSR_LOCK_WIDTH 1

/* REG_NSU_0_ING */
`define DDRMC5_NOC_REG_NSU_0_ING_OFFSET 17'h10
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ECC_CHK_EN 0
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ECC_CHK_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_DBI_EN 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_DBI_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOW_ORDER_EN 2
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOW_ORDER_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BEW_ORDER_EN 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BEW_ORDER_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_LLR_VC_MAP 6:4
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_LLR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED 7
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOR_VC_MAP 10:8
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_1 11
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BER_VC_MAP 14:12
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BER_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_2 15
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOW_VC_MAP 18:16
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_ISOW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_3 19
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BEW_VC_MAP 22:20
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_BEW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_4 31:23
`define DDRMC5_NOC_REG_NSU_0_ING_FLD_RESERVED_4_WIDTH 9
`define DDRMC5_NOC_REG_NSU_0_ING_WIDTH 23

/* REG_NSU_0_EGR */
`define DDRMC5_NOC_REG_NSU_0_EGR_OFFSET 17'h14
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_LLR_VC_MAP 2:0
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_LLR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISOR_VC_MAP 6:4
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISOR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_1 7
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BER_VC_MAP 10:8
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BER_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_2 11
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISOW_VC_MAP 14:12
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISOW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_3 15
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BEW_VC_MAP 18:16
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BEW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_4 19
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_4_WIDTH 1
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_LLR_PRI 21:20
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_LLR_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISR_PRI 23:22
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISR_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BER_PRI 25:24
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BER_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISW_PRI 27:26
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_ISW_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BEW_PRI 29:28
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_BEW_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_5 31:30
`define DDRMC5_NOC_REG_NSU_0_EGR_FLD_RESERVED_5_WIDTH 2
`define DDRMC5_NOC_REG_NSU_0_EGR_WIDTH 30

/* REG_NSU_1_ING */
`define DDRMC5_NOC_REG_NSU_1_ING_OFFSET 17'h18
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ECC_CHK_EN 0
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ECC_CHK_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_DBI_EN 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_DBI_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOW_ORDER_EN 2
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOW_ORDER_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BEW_ORDER_EN 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BEW_ORDER_EN_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_LLR_VC_MAP 6:4
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_LLR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED 7
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOR_VC_MAP 10:8
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_1 11
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BER_VC_MAP 14:12
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BER_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_2 15
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOW_VC_MAP 18:16
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_ISOW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_3 19
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BEW_VC_MAP 22:20
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_BEW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_4 31:23
`define DDRMC5_NOC_REG_NSU_1_ING_FLD_RESERVED_4_WIDTH 9
`define DDRMC5_NOC_REG_NSU_1_ING_WIDTH 23

/* REG_NSU_1_EGR */
`define DDRMC5_NOC_REG_NSU_1_EGR_OFFSET 17'h1c
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_LLR_VC_MAP 2:0
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_LLR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISOR_VC_MAP 6:4
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISOR_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_1 7
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_1_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BER_VC_MAP 10:8
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BER_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_2 11
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_2_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISOW_VC_MAP 14:12
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISOW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_3 15
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_3_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BEW_VC_MAP 18:16
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BEW_VC_MAP_WIDTH 3
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_4 19
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_4_WIDTH 1
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_LLR_PRI 21:20
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_LLR_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISR_PRI 23:22
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISR_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BER_PRI 25:24
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BER_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISW_PRI 27:26
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_ISW_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BEW_PRI 29:28
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_BEW_PRI_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_5 31:30
`define DDRMC5_NOC_REG_NSU_1_EGR_FLD_RESERVED_5_WIDTH 2
`define DDRMC5_NOC_REG_NSU_1_EGR_WIDTH 30

/* REG_TIMER_FIFO */
`define DDRMC5_NOC_REG_TIMER_FIFO_OFFSET 17'h20
`define DDRMC5_NOC_REG_TIMER_FIFO_FLD_DELAY_TAP 5:0
`define DDRMC5_NOC_REG_TIMER_FIFO_FLD_DELAY_TAP_WIDTH 6
`define DDRMC5_NOC_REG_TIMER_FIFO_FLD_RESERVED 31:6
`define DDRMC5_NOC_REG_TIMER_FIFO_FLD_RESERVED_WIDTH 26
`define DDRMC5_NOC_REG_TIMER_FIFO_WIDTH 6

/* REG_NSU0_PORT */
`define DDRMC5_NOC_REG_NSU0_PORT_OFFSET 17'h24
`define DDRMC5_NOC_REG_NSU0_PORT_FLD_SRC_ID 11:0
`define DDRMC5_NOC_REG_NSU0_PORT_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_REG_NSU0_PORT_FLD_RESERVED 31:12
`define DDRMC5_NOC_REG_NSU0_PORT_FLD_RESERVED_WIDTH 20
`define DDRMC5_NOC_REG_NSU0_PORT_WIDTH 12

/* REG_NSU1_PORT */
`define DDRMC5_NOC_REG_NSU1_PORT_OFFSET 17'h28
`define DDRMC5_NOC_REG_NSU1_PORT_FLD_SRC_ID 11:0
`define DDRMC5_NOC_REG_NSU1_PORT_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_REG_NSU1_PORT_FLD_RESERVED 31:12
`define DDRMC5_NOC_REG_NSU1_PORT_FLD_RESERVED_WIDTH 20
`define DDRMC5_NOC_REG_NSU1_PORT_WIDTH 12

/* REG_NSU_0_R_EGR */
`define DDRMC5_NOC_REG_NSU_0_R_EGR_OFFSET 17'h400
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_RESERVED 3:0
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_LLR_VC_TOKEN 11:4
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_LLR_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_ISOCR_VC_TOKEN 19:12
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_ISOCR_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_BER_VC_TOKEN 27:20
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_BER_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_RESERVED_1 31:28
`define DDRMC5_NOC_REG_NSU_0_R_EGR_FLD_RESERVED_1_WIDTH 4
`define DDRMC5_NOC_REG_NSU_0_R_EGR_WIDTH 28

/* REG_NSU_0_W_EGR */
`define DDRMC5_NOC_REG_NSU_0_W_EGR_OFFSET 17'h404
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_RESERVED 3:0
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_ISOCW_VC_TOKEN 11:4
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_ISOCW_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_BEW_VC_TOKEN 19:12
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_BEW_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_RESERVED_1 31:20
`define DDRMC5_NOC_REG_NSU_0_W_EGR_FLD_RESERVED_1_WIDTH 12
`define DDRMC5_NOC_REG_NSU_0_W_EGR_WIDTH 20

/* REG_NSU_1_R_EGR */
`define DDRMC5_NOC_REG_NSU_1_R_EGR_OFFSET 17'h408
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_RESERVED 3:0
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_LLR_VC_TOKEN 11:4
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_LLR_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_ISOCR_VC_TOKEN 19:12
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_ISOCR_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_BER_VC_TOKEN 27:20
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_BER_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_RESERVED_1 31:28
`define DDRMC5_NOC_REG_NSU_1_R_EGR_FLD_RESERVED_1_WIDTH 4
`define DDRMC5_NOC_REG_NSU_1_R_EGR_WIDTH 28

/* REG_NSU_1_W_EGR */
`define DDRMC5_NOC_REG_NSU_1_W_EGR_OFFSET 17'h40c
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_RESERVED 3:0
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_ISOCW_VC_TOKEN 11:4
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_ISOCW_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_BEW_VC_TOKEN 19:12
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_BEW_VC_TOKEN_WIDTH 8
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_RESERVED_1 31:20
`define DDRMC5_NOC_REG_NSU_1_W_EGR_FLD_RESERVED_1_WIDTH 12
`define DDRMC5_NOC_REG_NSU_1_W_EGR_WIDTH 20

/* REG_RD_DRR_TKN_P0 */
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_OFFSET 17'h410
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_LLR 7:0
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_LLR_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_ISOCR 15:8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_ISOCR_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_BER 23:16
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_BER_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_RESERVED 31:24
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_FLD_RESERVED_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P0_WIDTH 24

/* REG_WR_DRR_TKN_P0 */
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_OFFSET 17'h414
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_ISOCW 7:0
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_ISOCW_WIDTH 8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_BEW 15:8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_BEW_WIDTH 8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_RESERVED 31:16
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_REG_WR_DRR_TKN_P0_WIDTH 16

/* REG_RD_DRR_TKN_P1 */
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_OFFSET 17'h418
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_LLR 7:0
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_LLR_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_ISOCR 15:8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_ISOCR_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_BER 23:16
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_BER_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_RESERVED 31:24
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_FLD_RESERVED_WIDTH 8
`define DDRMC5_NOC_REG_RD_DRR_TKN_P1_WIDTH 24

/* REG_WR_DRR_TKN_P1 */
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_OFFSET 17'h41c
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_ISOCW 7:0
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_ISOCW_WIDTH 8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_BEW 15:8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_BEW_WIDTH 8
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_RESERVED 31:16
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_REG_WR_DRR_TKN_P1_WIDTH 16

/* REG_QOS0 */
`define DDRMC5_NOC_REG_QOS0_OFFSET 17'h420
`define DDRMC5_NOC_REG_QOS0_FLD_ARB_MODE 0
`define DDRMC5_NOC_REG_QOS0_FLD_ARB_MODE_WIDTH 1
`define DDRMC5_NOC_REG_QOS0_FLD_RESERVED 3:1
`define DDRMC5_NOC_REG_QOS0_FLD_RESERVED_WIDTH 3
`define DDRMC5_NOC_REG_QOS0_FLD_RD_THRSHOLD 15:4
`define DDRMC5_NOC_REG_QOS0_FLD_RD_THRSHOLD_WIDTH 12
`define DDRMC5_NOC_REG_QOS0_FLD_WR_THRSHOLD 27:16
`define DDRMC5_NOC_REG_QOS0_FLD_WR_THRSHOLD_WIDTH 12
`define DDRMC5_NOC_REG_QOS0_FLD_RESERVED_1 31:28
`define DDRMC5_NOC_REG_QOS0_FLD_RESERVED_1_WIDTH 4
`define DDRMC5_NOC_REG_QOS0_WIDTH 28

/* REG_QOS1 */
`define DDRMC5_NOC_REG_QOS1_OFFSET 17'h424
`define DDRMC5_NOC_REG_QOS1_FLD_LLR_TOKEN 9:0
`define DDRMC5_NOC_REG_QOS1_FLD_LLR_TOKEN_WIDTH 10
`define DDRMC5_NOC_REG_QOS1_FLD_ISOR_TOKEN 19:10
`define DDRMC5_NOC_REG_QOS1_FLD_ISOR_TOKEN_WIDTH 10
`define DDRMC5_NOC_REG_QOS1_FLD_BER_TOKEN 29:20
`define DDRMC5_NOC_REG_QOS1_FLD_BER_TOKEN_WIDTH 10
`define DDRMC5_NOC_REG_QOS1_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_QOS1_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_QOS1_WIDTH 30

/* REG_QOS2 */
`define DDRMC5_NOC_REG_QOS2_OFFSET 17'h428
`define DDRMC5_NOC_REG_QOS2_FLD_ISOW_TOKEN 9:0
`define DDRMC5_NOC_REG_QOS2_FLD_ISOW_TOKEN_WIDTH 10
`define DDRMC5_NOC_REG_QOS2_FLD_BEW_TOKEN 19:10
`define DDRMC5_NOC_REG_QOS2_FLD_BEW_TOKEN_WIDTH 10
`define DDRMC5_NOC_REG_QOS2_FLD_RESERVED 31:20
`define DDRMC5_NOC_REG_QOS2_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_REG_QOS2_WIDTH 20

/* REG_QOS_TIMEOUT0 */
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_OFFSET 17'h42c
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_LLR_SCALE 4:0
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_LLR_SCALE_WIDTH 5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_ISR_SCALE 9:5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_ISR_SCALE_WIDTH 5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_BER_SCALE 14:10
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_BER_SCALE_WIDTH 5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_ISW_SCALE 19:15
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_ISW_SCALE_WIDTH 5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_BEW_SCALE 24:20
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_BEW_SCALE_WIDTH 5
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_RESERVED 31:25
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_REG_QOS_TIMEOUT0_WIDTH 25

/* REG_QOS_TIMEOUT1 */
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_OFFSET 17'h430
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_LLR_TIMEOUT 7:0
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_LLR_TIMEOUT_WIDTH 8
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_ISOR_TIMEOUT 15:8
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_ISOR_TIMEOUT_WIDTH 8
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_BER_TIMEOUT 23:16
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_BER_TIMEOUT_WIDTH 8
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_ISOW_TIMEOUT 31:24
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_FLD_ISOW_TIMEOUT_WIDTH 8
`define DDRMC5_NOC_REG_QOS_TIMEOUT1_WIDTH 32

/* REG_QOS_TIMEOUT2 */
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_OFFSET 17'h434
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_FLD_BEW_TIMEOUT 7:0
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_FLD_BEW_TIMEOUT_WIDTH 8
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_FLD_RESERVED 31:8
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_FLD_RESERVED_WIDTH 24
`define DDRMC5_NOC_REG_QOS_TIMEOUT2_WIDTH 8

/* REG_RATE_CTRL_SCALE */
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_OFFSET 17'h438
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_LLR_UPDATE_PERIOD 4:0
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_LLR_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_ISR_UPDATE_PERIOD 9:5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_ISR_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_BER_UPDATE_PERIOD 14:10
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_BER_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_ISW_UPDATE_PERIOD 19:15
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_ISW_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_BEW_UPDATE_PERIOD 24:20
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_BEW_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_RESERVED 31:25
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_REG_RATE_CTRL_SCALE_WIDTH 25

/* REG_P0_LLR_RATE_CTRL */
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_OFFSET 17'h43c
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P0_LLR_RATE_CTRL_WIDTH 22

/* REG_P0_ISR_RATE_CTRL */
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_OFFSET 17'h440
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P0_ISR_RATE_CTRL_WIDTH 22

/* REG_P0_BER_RATE_CTRL */
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_OFFSET 17'h444
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P0_BER_RATE_CTRL_WIDTH 22

/* REG_P0_ISW_RATE_CTRL */
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_OFFSET 17'h448
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P0_ISW_RATE_CTRL_WIDTH 22

/* REG_P0_BEW_RATE_CTRL */
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_OFFSET 17'h44c
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P0_BEW_RATE_CTRL_WIDTH 22

/* REG_P1_LLR_RATE_CTRL */
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_OFFSET 17'h450
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P1_LLR_RATE_CTRL_WIDTH 22

/* REG_P1_ISR_RATE_CTRL */
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_OFFSET 17'h454
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P1_ISR_RATE_CTRL_WIDTH 22

/* REG_P1_BER_RATE_CTRL */
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_OFFSET 17'h458
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P1_BER_RATE_CTRL_WIDTH 22

/* REG_P1_ISW_RATE_CTRL */
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_OFFSET 17'h45c
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P1_ISW_RATE_CTRL_WIDTH 22

/* REG_P1_BEW_RATE_CTRL */
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_OFFSET 17'h460
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_P1_BEW_RATE_CTRL_WIDTH 22

/* REG_SCRUB_WAIT */
`define DDRMC5_NOC_REG_SCRUB_WAIT_OFFSET 17'h464
`define DDRMC5_NOC_REG_SCRUB_WAIT_FLD_CNT 7:0
`define DDRMC5_NOC_REG_SCRUB_WAIT_FLD_CNT_WIDTH 8
`define DDRMC5_NOC_REG_SCRUB_WAIT_FLD_RESERVED 31:8
`define DDRMC5_NOC_REG_SCRUB_WAIT_FLD_RESERVED_WIDTH 24
`define DDRMC5_NOC_REG_SCRUB_WAIT_WIDTH 8

/* REG_CMDQ_LLR_RATE_CTRL */
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_OFFSET 17'h468
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_LLR_RATE_CTRL_WIDTH 22

/* REG_CMDQ_ISR_RATE_CTRL */
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_OFFSET 17'h46c
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_ISR_RATE_CTRL_WIDTH 22

/* REG_CMDQ_BER_RATE_CTRL */
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_OFFSET 17'h470
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_BER_RATE_CTRL_WIDTH 22

/* REG_CMDQ_ISW_RATE_CTRL */
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_OFFSET 17'h474
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_ISW_RATE_CTRL_WIDTH 22

/* REG_CMDQ_BEW_RATE_CTRL */
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_OFFSET 17'h478
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_CREDIT_UPDATE 9:0
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_CREDIT_UPDATE_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_CREDIT_LIMIT 21:10
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_CREDIT_LIMIT_WIDTH 12
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_RESERVED 31:22
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_CMDQ_BEW_RATE_CTRL_WIDTH 22

/* REG_QOS_RATE_CTRL_SCALE */
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_OFFSET 17'h47c
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_LLR_UPDATE_PERIOD 4:0
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_LLR_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_ISR_UPDATE_PERIOD 9:5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_ISR_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_BER_UPDATE_PERIOD 14:10
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_BER_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_ISW_UPDATE_PERIOD 19:15
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_ISW_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_BEW_UPDATE_PERIOD 24:20
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_BEW_UPDATE_PERIOD_WIDTH 5
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_RESERVED 31:25
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_REG_QOS_RATE_CTRL_SCALE_WIDTH 25

/* EXMON_CLR_EXE */
`define DDRMC5_NOC_EXMON_CLR_EXE_OFFSET 17'h480
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_0 0
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_0_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_1 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_1_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_2 2
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_2_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_3 3
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_3_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_4 4
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_4_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_5 5
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_5_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_6 6
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_6_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_7 7
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_MON_7_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_AXSIZE_BASED_CHECK 8
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_AXSIZE_BASED_CHECK_WIDTH 1
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_RESERVED 31:9
`define DDRMC5_NOC_EXMON_CLR_EXE_FLD_RESERVED_WIDTH 23
`define DDRMC5_NOC_EXMON_CLR_EXE_WIDTH 9

/* UB_CLK_MUX */
`define DDRMC5_NOC_UB_CLK_MUX_OFFSET 17'h484
`define DDRMC5_NOC_UB_CLK_MUX_FLD_SEL 1:0
`define DDRMC5_NOC_UB_CLK_MUX_FLD_SEL_WIDTH 2
`define DDRMC5_NOC_UB_CLK_MUX_FLD_RESERVED 31:2
`define DDRMC5_NOC_UB_CLK_MUX_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_UB_CLK_MUX_WIDTH 2

/* NSU0_PERF_MON_CTL_0_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_OFFSET 17'h488
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_MON_EN 0
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_MON_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_SNGL 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_SNGL_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_RESERVED 31:2
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_0_WIDTH 2

/* NSU0_PERF_MON_CTL_0_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_OFFSET 17'h48c
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_TB_SEL 2:0
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_TB_SEL_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_LAT_SEL 3
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_LAT_SEL_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_LLR 4
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_LLR_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_ISOR 5
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_ISOR_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_BER 6
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_BER_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_ISOW 7
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_ISOW_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_BEW 8
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_BEW_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_RESERVED 31:9
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_FLD_RESERVED_WIDTH 23
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_0_1_WIDTH 9

/* NSU0_PERF_FILTER_0_0 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_OFFSET 17'h490
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXID 15:0
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXID_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLEN_MIN 19:16
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLEN_MIN_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLEN_MAX 23:20
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLEN_MAX_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXBURST 25:24
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXPROT 28:26
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXPROT_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLOCK 29
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_RESERVED 31:30
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_0_WIDTH 30

/* NSU0_PERF_FILTER_0_1 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_OFFSET 17'h494
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_SRC_ID 11:0
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_SMID 21:12
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_RESERVED 31:22
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_NSU0_PERF_FILTER_0_1_WIDTH 22

/* NSU0_PERF_FILTER_EN_0 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_OFFSET 17'h498
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXID 0
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXLEN 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXLEN_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXBURST 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXBURST_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXPROT 3
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXPROT_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXLOCK 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_SRC_ID 5
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_SRC_ID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_SMID 6
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_SMID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_RESERVED 31:7
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_0_WIDTH 7

/* NSU0_PERF_MON_0_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_0_OFFSET 17'h49c
`define DDRMC5_NOC_NSU0_PERF_MON_0_0_FLD_LAT_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_0_FLD_LAT_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_0_0_WIDTH 32

/* NSU0_PERF_MON_0_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_OFFSET 17'h4a0
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_LAT_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_LAT_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_LAT_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_LAT_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_0_1_WIDTH 17

/* NSU0_PERF_MON_0_2 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_2_OFFSET 17'h4a4
`define DDRMC5_NOC_NSU0_PERF_MON_0_2_FLD_BURST_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_2_FLD_BURST_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_0_2_WIDTH 32

/* NSU0_PERF_MON_0_3 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_OFFSET 17'h4a8
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_FLD_BURST_HI 30:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_FLD_BURST_HI_WIDTH 31
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_FLD_BURST_OVF 31
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_FLD_BURST_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_0_3_WIDTH 32

/* NSU0_PERF_MON_0_4 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_4_OFFSET 17'h4ac
`define DDRMC5_NOC_NSU0_PERF_MON_0_4_FLD_HEADER_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_4_FLD_HEADER_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_0_4_WIDTH 32

/* NSU0_PERF_MON_0_5 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_OFFSET 17'h4b0
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_HEADER_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_HEADER_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_HEADER_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_HEADER_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_0_5_WIDTH 17

/* NSU0_PERF_MON_0_ROLLOVER */
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_OFFSET 17'h4b4
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_FLD_CURNT_TIME_ROLLOVER 3:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_FLD_CURNT_TIME_ROLLOVER_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_FLD_RESERVED 31:4
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_NSU0_PERF_MON_0_ROLLOVER_WIDTH 4

/* NSU0_PERF_MON_0_START_TIME_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_0_OFFSET 17'h4b8
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_0_WIDTH 32

/* NSU0_PERF_MON_0_START_TIME_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_OFFSET 17'h4bc
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_FLD_INTERVAL_TIME_HI 2:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_FLD_RESERVED 31:3
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_FLD_RESERVED_WIDTH 29
`define DDRMC5_NOC_NSU0_PERF_MON_0_START_TIME_1_WIDTH 3

/* NSU0_PERF_MON_0_STOP_TIME_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_0_OFFSET 17'h4c0
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_0_WIDTH 32

/* NSU0_PERF_MON_0_STOP_TIME_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_OFFSET 17'h4c4
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_0_STOP_TIME_1_WIDTH 17

/* NSU0_PERF_MON_CTL_1_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_OFFSET 17'h4c8
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_MON_EN 0
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_MON_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_SNGL 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_SNGL_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_RESERVED 31:2
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_0_WIDTH 2

/* NSU0_PERF_MON_CTL_1_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_OFFSET 17'h4cc
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_TB_SEL 2:0
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_TB_SEL_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_LAT_SEL 3
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_LAT_SEL_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_LLR 4
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_LLR_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_ISOR 5
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_ISOR_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_BER 6
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_BER_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_ISOW 7
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_ISOW_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_BEW 8
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_BEW_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_RESERVED 31:9
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_FLD_RESERVED_WIDTH 23
`define DDRMC5_NOC_NSU0_PERF_MON_CTL_1_1_WIDTH 9

/* NSU0_PERF_FILTER_1_0 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_OFFSET 17'h4d0
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXID 15:0
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXID_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLEN_MIN 19:16
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLEN_MIN_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLEN_MAX 23:20
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLEN_MAX_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXBURST 25:24
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXPROT 28:26
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXPROT_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLOCK 29
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_RESERVED 31:30
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_0_WIDTH 30

/* NSU0_PERF_FILTER_1_1 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_OFFSET 17'h4d4
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_SRC_ID 11:0
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_SMID 21:12
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_RESERVED 31:22
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_NSU0_PERF_FILTER_1_1_WIDTH 22

/* NSU0_PERF_FILTER_EN_1 */
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_OFFSET 17'h4d8
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXID 0
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXLEN 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXLEN_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXBURST 2
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXBURST_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXPROT 3
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXPROT_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXLOCK 4
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_SRC_ID 5
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_SRC_ID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_SMID 6
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_SMID_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_RESERVED 31:7
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_NSU0_PERF_FILTER_EN_1_WIDTH 7

/* NSU0_PERF_MON_1_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_0_OFFSET 17'h4dc
`define DDRMC5_NOC_NSU0_PERF_MON_1_0_FLD_LAT_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_0_FLD_LAT_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_1_0_WIDTH 32

/* NSU0_PERF_MON_1_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_OFFSET 17'h4e0
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_LAT_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_LAT_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_LAT_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_LAT_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_1_1_WIDTH 17

/* NSU0_PERF_MON_1_2 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_2_OFFSET 17'h4e4
`define DDRMC5_NOC_NSU0_PERF_MON_1_2_FLD_BURST_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_2_FLD_BURST_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_1_2_WIDTH 32

/* NSU0_PERF_MON_1_3 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_OFFSET 17'h4e8
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_FLD_BURST_HI 30:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_FLD_BURST_HI_WIDTH 31
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_FLD_BURST_OVF 31
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_FLD_BURST_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_1_3_WIDTH 32

/* NSU0_PERF_MON_1_4 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_4_OFFSET 17'h4ec
`define DDRMC5_NOC_NSU0_PERF_MON_1_4_FLD_HEADER_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_4_FLD_HEADER_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_1_4_WIDTH 32

/* NSU0_PERF_MON_1_5 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_OFFSET 17'h4f0
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_HEADER_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_HEADER_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_HEADER_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_HEADER_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_1_5_WIDTH 17

/* NSU0_PERF_MON_1_ROLLOVER */
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_OFFSET 17'h4f4
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_FLD_CURNT_TIME_ROLLOVER 3:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_FLD_CURNT_TIME_ROLLOVER_WIDTH 4
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_FLD_RESERVED 31:4
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_NSU0_PERF_MON_1_ROLLOVER_WIDTH 4

/* NSU0_PERF_MON_1_START_TIME_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_0_OFFSET 17'h4f8
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_0_WIDTH 32

/* NSU0_PERF_MON_1_START_TIME_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_OFFSET 17'h4fc
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_FLD_INTERVAL_TIME_HI 2:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 3
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_FLD_RESERVED 31:3
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_FLD_RESERVED_WIDTH 29
`define DDRMC5_NOC_NSU0_PERF_MON_1_START_TIME_1_WIDTH 3

/* NSU0_PERF_MON_1_STOP_TIME_0 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_0_OFFSET 17'h500
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_0_WIDTH 32

/* NSU0_PERF_MON_1_STOP_TIME_1 */
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_OFFSET 17'h504
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI 15:0
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF 16
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF_WIDTH 1
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU0_PERF_MON_1_STOP_TIME_1_WIDTH 17

/* NSU1_PERF_MON_CTL_0_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_OFFSET 17'h508
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_MON_EN 0
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_MON_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_SNGL 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_SNGL_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_RESERVED 31:2
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_0_WIDTH 2

/* NSU1_PERF_MON_CTL_0_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_OFFSET 17'h50c
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_TB_SEL 2:0
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_TB_SEL_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_LAT_SEL 3
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_LAT_SEL_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_LLR 4
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_LLR_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_ISOR 5
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_ISOR_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_BER 6
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_BER_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_ISOW 7
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_ISOW_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_BEW 8
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_BEW_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_RESERVED 31:9
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_FLD_RESERVED_WIDTH 23
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_0_1_WIDTH 9

/* NSU1_PERF_FILTER_0_0 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_OFFSET 17'h510
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXID 15:0
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXID_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLEN_MIN 19:16
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLEN_MIN_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLEN_MAX 23:20
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLEN_MAX_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXBURST 25:24
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXPROT 28:26
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXPROT_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLOCK 29
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_RESERVED 31:30
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_0_WIDTH 30

/* NSU1_PERF_FILTER_0_1 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_OFFSET 17'h514
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_SRC_ID 11:0
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_SMID 21:12
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_RESERVED 31:22
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_NSU1_PERF_FILTER_0_1_WIDTH 22

/* NSU1_PERF_FILTER_EN_0 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_OFFSET 17'h518
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXID 0
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXLEN 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXLEN_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXBURST 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXBURST_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXPROT 3
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXPROT_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXLOCK 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_SRC_ID 5
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_SRC_ID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_SMID 6
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_SMID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_RESERVED 31:7
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_0_WIDTH 7

/* NSU1_PERF_MON_0_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_0_OFFSET 17'h51c
`define DDRMC5_NOC_NSU1_PERF_MON_0_0_FLD_LAT_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_0_FLD_LAT_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_0_0_WIDTH 32

/* NSU1_PERF_MON_0_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_OFFSET 17'h520
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_LAT_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_LAT_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_LAT_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_LAT_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_0_1_WIDTH 17

/* NSU1_PERF_MON_0_2 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_2_OFFSET 17'h524
`define DDRMC5_NOC_NSU1_PERF_MON_0_2_FLD_BURST_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_2_FLD_BURST_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_0_2_WIDTH 32

/* NSU1_PERF_MON_0_3 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_OFFSET 17'h528
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_FLD_BURST_HI 30:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_FLD_BURST_HI_WIDTH 31
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_FLD_BURST_OVF 31
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_FLD_BURST_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_0_3_WIDTH 32

/* NSU1_PERF_MON_0_4 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_4_OFFSET 17'h52c
`define DDRMC5_NOC_NSU1_PERF_MON_0_4_FLD_HEADER_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_4_FLD_HEADER_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_0_4_WIDTH 32

/* NSU1_PERF_MON_0_5 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_OFFSET 17'h530
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_HEADER_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_HEADER_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_HEADER_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_HEADER_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_0_5_WIDTH 17

/* NSU1_PERF_MON_0_ROLLOVER */
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_OFFSET 17'h534
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_FLD_CURNT_TIME_ROLLOVER 3:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_FLD_CURNT_TIME_ROLLOVER_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_FLD_RESERVED 31:4
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_NSU1_PERF_MON_0_ROLLOVER_WIDTH 4

/* NSU1_PERF_MON_0_START_TIME_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_0_OFFSET 17'h538
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_0_WIDTH 32

/* NSU1_PERF_MON_0_START_TIME_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_OFFSET 17'h53c
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_FLD_INTERVAL_TIME_HI 2:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_FLD_RESERVED 31:3
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_FLD_RESERVED_WIDTH 29
`define DDRMC5_NOC_NSU1_PERF_MON_0_START_TIME_1_WIDTH 3

/* NSU1_PERF_MON_0_STOP_TIME_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_0_OFFSET 17'h540
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_0_WIDTH 32

/* NSU1_PERF_MON_0_STOP_TIME_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_OFFSET 17'h544
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_0_STOP_TIME_1_WIDTH 17

/* NSU1_PERF_MON_CTL_1_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_OFFSET 17'h548
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_MON_EN 0
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_MON_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_SNGL 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_SNGL_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_RESERVED 31:2
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_0_WIDTH 2

/* NSU1_PERF_MON_CTL_1_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_OFFSET 17'h54c
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_TB_SEL 2:0
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_TB_SEL_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_LAT_SEL 3
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_LAT_SEL_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_LLR 4
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_LLR_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_ISOR 5
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_ISOR_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_BER 6
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_BER_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_ISOW 7
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_ISOW_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_BEW 8
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_BEW_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_RESERVED 31:9
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_FLD_RESERVED_WIDTH 23
`define DDRMC5_NOC_NSU1_PERF_MON_CTL_1_1_WIDTH 9

/* NSU1_PERF_FILTER_1_0 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_OFFSET 17'h550
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXID 15:0
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXID_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLEN_MIN 19:16
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLEN_MIN_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLEN_MAX 23:20
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLEN_MAX_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXBURST 25:24
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXPROT 28:26
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXPROT_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLOCK 29
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_RESERVED 31:30
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_0_WIDTH 30

/* NSU1_PERF_FILTER_1_1 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_OFFSET 17'h554
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_SRC_ID 11:0
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_SRC_ID_WIDTH 12
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_SMID 21:12
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_RESERVED 31:22
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_NSU1_PERF_FILTER_1_1_WIDTH 22

/* NSU1_PERF_FILTER_EN_1 */
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_OFFSET 17'h558
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXID 0
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXLEN 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXLEN_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXBURST 2
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXBURST_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXPROT 3
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXPROT_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXLOCK 4
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_SRC_ID 5
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_SRC_ID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_SMID 6
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_SMID_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_RESERVED 31:7
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_NSU1_PERF_FILTER_EN_1_WIDTH 7

/* NSU1_PERF_MON_1_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_0_OFFSET 17'h55c
`define DDRMC5_NOC_NSU1_PERF_MON_1_0_FLD_LAT_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_0_FLD_LAT_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_1_0_WIDTH 32

/* NSU1_PERF_MON_1_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_OFFSET 17'h560
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_LAT_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_LAT_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_LAT_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_LAT_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_1_1_WIDTH 17

/* NSU1_PERF_MON_1_2 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_2_OFFSET 17'h564
`define DDRMC5_NOC_NSU1_PERF_MON_1_2_FLD_BURST_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_2_FLD_BURST_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_1_2_WIDTH 32

/* NSU1_PERF_MON_1_3 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_OFFSET 17'h568
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_FLD_BURST_HI 30:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_FLD_BURST_HI_WIDTH 31
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_FLD_BURST_OVF 31
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_FLD_BURST_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_1_3_WIDTH 32

/* NSU1_PERF_MON_1_4 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_4_OFFSET 17'h56c
`define DDRMC5_NOC_NSU1_PERF_MON_1_4_FLD_HEADER_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_4_FLD_HEADER_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_1_4_WIDTH 32

/* NSU1_PERF_MON_1_5 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_OFFSET 17'h570
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_HEADER_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_HEADER_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_HEADER_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_HEADER_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_1_5_WIDTH 17

/* NSU1_PERF_MON_1_ROLLOVER */
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_OFFSET 17'h574
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_FLD_CURNT_TIME_ROLLOVER 3:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_FLD_CURNT_TIME_ROLLOVER_WIDTH 4
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_FLD_RESERVED 31:4
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_NSU1_PERF_MON_1_ROLLOVER_WIDTH 4

/* NSU1_PERF_MON_1_START_TIME_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_0_OFFSET 17'h578
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_0_WIDTH 32

/* NSU1_PERF_MON_1_START_TIME_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_OFFSET 17'h57c
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_FLD_INTERVAL_TIME_HI 2:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 3
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_FLD_RESERVED 31:3
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_FLD_RESERVED_WIDTH 29
`define DDRMC5_NOC_NSU1_PERF_MON_1_START_TIME_1_WIDTH 3

/* NSU1_PERF_MON_1_STOP_TIME_0 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_0_OFFSET 17'h580
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_0_FLD_INTERVAL_TIME_LOW 31:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_0_FLD_INTERVAL_TIME_LOW_WIDTH 32
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_0_WIDTH 32

/* NSU1_PERF_MON_1_STOP_TIME_1 */
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_OFFSET 17'h584
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI 15:0
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_WIDTH 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF 16
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_INTERVAL_TIME_HI_OVF_WIDTH 1
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_RESERVED 31:17
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_FLD_RESERVED_WIDTH 15
`define DDRMC5_NOC_NSU1_PERF_MON_1_STOP_TIME_1_WIDTH 17

/* NSU0_ERR_LOG0_EN */
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_OFFSET 17'h588
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_ING_OF 12
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU0_ERR_LOG0_EN_WIDTH 25

/* NSU0_ERR_LOG1_EN */
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_OFFSET 17'h58c
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_ING_OF 12
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU0_ERR_LOG1_EN_WIDTH 25

/* NSU0_ERR_STATUS */
`define DDRMC5_NOC_NSU0_ERR_STATUS_OFFSET 17'h590
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_ING_OF 12
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU0_ERR_STATUS_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU0_ERR_STATUS_WIDTH 25

/* NSU0_ERR_LOG0_0 */
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_OFFSET 17'h594
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_TAG 7:0
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_TAG_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_SRC 19:8
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_SRC_WIDTH 12
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_DST 31:20
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_FLD_DST_WIDTH 12
`define DDRMC5_NOC_NSU0_ERR_LOG0_0_WIDTH 32

/* NSU0_ERR_LOG0_1 */
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_OFFSET 17'h598
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_PKT_TYPE 3:0
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_PKT_TYPE_WIDTH 4
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_DST_PAR 4
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_DST_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_WSTRB 20:5
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_WSTRB_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_LAST 21
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_LAST_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_VC 26:22
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_VC_WIDTH 5
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_RESERVED 30:27
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_POISON 31
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_FLD_POISON_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_1_WIDTH 32

/* NSU0_ERR_LOG0_2 */
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_OFFSET 17'h59c
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_NPP_EBIT 7:0
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_NPP_EBIT_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXLEN 15:8
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXLEN_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXSIZE 18:16
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXSIZE_WIDTH 3
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXLOCK 19
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_SMID 29:20
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXBURST 31:30
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU0_ERR_LOG0_2_WIDTH 32

/* NSU0_ERR_LOG0_3 */
`define DDRMC5_NOC_NSU0_ERR_LOG0_3_OFFSET 17'h5a0
`define DDRMC5_NOC_NSU0_ERR_LOG0_3_FLD_ADDR_L 31:0
`define DDRMC5_NOC_NSU0_ERR_LOG0_3_FLD_ADDR_L_WIDTH 32
`define DDRMC5_NOC_NSU0_ERR_LOG0_3_WIDTH 32

/* NSU0_ERR_LOG0_4 */
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_OFFSET 17'h5a4
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_FLD_ADDR_U 15:0
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_FLD_ADDR_U_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_FLD_ERR_REF_NUM 31:16
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_FLD_ERR_REF_NUM_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG0_4_WIDTH 32

/* NSU0_ERR_LOG1_0 */
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_OFFSET 17'h5a8
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_TAG 7:0
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_TAG_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_SRC 19:8
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_SRC_WIDTH 12
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_DST 31:20
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_FLD_DST_WIDTH 12
`define DDRMC5_NOC_NSU0_ERR_LOG1_0_WIDTH 32

/* NSU0_ERR_LOG1_1 */
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_OFFSET 17'h5ac
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_PKT_TYPE 3:0
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_PKT_TYPE_WIDTH 4
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_DST_PAR 4
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_DST_PAR_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_WSTRB 20:5
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_WSTRB_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_LAST 21
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_LAST_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_VC 26:22
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_VC_WIDTH 5
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_RESERVED 30:27
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_POISON 31
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_FLD_POISON_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_1_WIDTH 32

/* NSU0_ERR_LOG1_2 */
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_OFFSET 17'h5b0
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_NPP_EBIT 7:0
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_NPP_EBIT_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXLEN 15:8
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXLEN_WIDTH 8
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXSIZE 18:16
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXSIZE_WIDTH 3
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXLOCK 19
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_SMID 29:20
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXBURST 31:30
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU0_ERR_LOG1_2_WIDTH 32

/* NSU0_ERR_LOG1_3 */
`define DDRMC5_NOC_NSU0_ERR_LOG1_3_OFFSET 17'h5b4
`define DDRMC5_NOC_NSU0_ERR_LOG1_3_FLD_ADDR_L 31:0
`define DDRMC5_NOC_NSU0_ERR_LOG1_3_FLD_ADDR_L_WIDTH 32
`define DDRMC5_NOC_NSU0_ERR_LOG1_3_WIDTH 32

/* NSU0_ERR_LOG1_4 */
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_OFFSET 17'h5b8
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_FLD_ADDR_U 15:0
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_FLD_ADDR_U_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_FLD_ERR_REF_NUM 31:16
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_FLD_ERR_REF_NUM_WIDTH 16
`define DDRMC5_NOC_NSU0_ERR_LOG1_4_WIDTH 32

/* NSU1_ERR_LOG0_EN */
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_OFFSET 17'h5bc
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_ING_OF 12
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU1_ERR_LOG0_EN_WIDTH 25

/* NSU1_ERR_LOG1_EN */
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_OFFSET 17'h5c0
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_ING_OF 12
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU1_ERR_LOG1_EN_WIDTH 25

/* NSU1_ERR_STATUS */
`define DDRMC5_NOC_NSU1_ERR_STATUS_OFFSET 17'h5c4
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_UNALIGN_WRAP 0
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_UNALIGN_WRAP_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_SIZE_INVALID 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EX_SIZE_INVALID 2
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EX_SIZE_INVALID_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_WRAP_LEN 3
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_WRAP_LEN 4
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_WRAP_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_DBI_ID_PAR 5
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_DBI_ID_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_UC 6
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_UC 7
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_UNMAP_VC 8
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_UNMAP_VC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_DST_ID_MATCH 9
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_DST_ID_MATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_NUM_LEN 10
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_NUM_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EGR_OF 11
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EGR_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_ING_OF 12
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_ING_OF_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EX_LEN 13
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_EX_LEN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_RESP_PAR 14
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_RESP_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_UC 15
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_UC_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_CE 16
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_CE 17
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_CE 18
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_2ND_CE 19
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_2ND_CE 20
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_2ND_CE 21
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RD_HEADER_2ND_CE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_POISON 22
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_WR_DATA_POISON_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_VC_TYP_MISSMATCH 23
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_VC_TYP_MISSMATCH_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_NOT_READY 24
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_NOT_READY_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RESERVED 31:25
`define DDRMC5_NOC_NSU1_ERR_STATUS_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_NSU1_ERR_STATUS_WIDTH 25

/* NSU1_ERR_LOG0_0 */
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_OFFSET 17'h5c8
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_TAG 7:0
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_TAG_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_SRC 19:8
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_SRC_WIDTH 12
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_DST 31:20
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_FLD_DST_WIDTH 12
`define DDRMC5_NOC_NSU1_ERR_LOG0_0_WIDTH 32

/* NSU1_ERR_LOG0_1 */
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_OFFSET 17'h5cc
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_PKT_TYPE 3:0
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_PKT_TYPE_WIDTH 4
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_DST_PAR 4
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_DST_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_WSTRB 20:5
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_WSTRB_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_LAST 21
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_LAST_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_VC 26:22
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_VC_WIDTH 5
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_RESERVED 30:27
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_POISON 31
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_FLD_POISON_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_1_WIDTH 32

/* NSU1_ERR_LOG0_2 */
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_OFFSET 17'h5d0
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_NPP_EBIT 7:0
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_NPP_EBIT_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXLEN 15:8
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXLEN_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXSIZE 18:16
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXSIZE_WIDTH 3
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXLOCK 19
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_SMID 29:20
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXBURST 31:30
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU1_ERR_LOG0_2_WIDTH 32

/* NSU1_ERR_LOG0_3 */
`define DDRMC5_NOC_NSU1_ERR_LOG0_3_OFFSET 17'h5d4
`define DDRMC5_NOC_NSU1_ERR_LOG0_3_FLD_ADDR_L 31:0
`define DDRMC5_NOC_NSU1_ERR_LOG0_3_FLD_ADDR_L_WIDTH 32
`define DDRMC5_NOC_NSU1_ERR_LOG0_3_WIDTH 32

/* NSU1_ERR_LOG0_4 */
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_OFFSET 17'h5d8
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_FLD_ADDR_U 15:0
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_FLD_ADDR_U_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_FLD_ERR_REF_NUM 31:16
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_FLD_ERR_REF_NUM_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG0_4_WIDTH 32

/* NSU1_ERR_LOG1_0 */
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_OFFSET 17'h5dc
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_TAG 7:0
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_TAG_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_SRC 19:8
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_SRC_WIDTH 12
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_DST 31:20
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_FLD_DST_WIDTH 12
`define DDRMC5_NOC_NSU1_ERR_LOG1_0_WIDTH 32

/* NSU1_ERR_LOG1_1 */
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_OFFSET 17'h5e0
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_PKT_TYPE 3:0
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_PKT_TYPE_WIDTH 4
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_DST_PAR 4
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_DST_PAR_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_WSTRB 20:5
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_WSTRB_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_LAST 21
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_LAST_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_VC 26:22
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_VC_WIDTH 5
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_RESERVED 30:27
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_POISON 31
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_FLD_POISON_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_1_WIDTH 32

/* NSU1_ERR_LOG1_2 */
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_OFFSET 17'h5e4
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_NPP_EBIT 7:0
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_NPP_EBIT_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXLEN 15:8
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXLEN_WIDTH 8
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXSIZE 18:16
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXSIZE_WIDTH 3
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXLOCK 19
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXLOCK_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_SMID 29:20
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_SMID_WIDTH 10
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXBURST 31:30
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_FLD_AXBURST_WIDTH 2
`define DDRMC5_NOC_NSU1_ERR_LOG1_2_WIDTH 32

/* NSU1_ERR_LOG1_3 */
`define DDRMC5_NOC_NSU1_ERR_LOG1_3_OFFSET 17'h5e8
`define DDRMC5_NOC_NSU1_ERR_LOG1_3_FLD_ADDR_L 31:0
`define DDRMC5_NOC_NSU1_ERR_LOG1_3_FLD_ADDR_L_WIDTH 32
`define DDRMC5_NOC_NSU1_ERR_LOG1_3_WIDTH 32

/* NSU1_ERR_LOG1_4 */
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_OFFSET 17'h5ec
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_FLD_ADDR_U 15:0
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_FLD_ADDR_U_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_FLD_ERR_REF_NUM 31:16
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_FLD_ERR_REF_NUM_WIDTH 16
`define DDRMC5_NOC_NSU1_ERR_LOG1_4_WIDTH 32

/* NSU0_ERR_CTRL */
`define DDRMC5_NOC_NSU0_ERR_CTRL_OFFSET 17'h5f0
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_RESERVED 11:0
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_PAR_RESP_ERR_EN 12
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_PAR_RESP_ERR_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_FATAL_DROP_EN 13
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_FATAL_DROP_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_SEL 15:14
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_SEL_WIDTH 2
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_DW_EN 16
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_DW_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_CW_EN 17
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_CW_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_R_EN 18
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_R_EN_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_DW_DONE 19
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_DW_DONE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_CW_DONE 20
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_CW_DONE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_R_DONE 21
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_R_DONE_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_PERSISTENT 22
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_PERSISTENT_WIDTH 1
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_RESERVED_1 31:23
`define DDRMC5_NOC_NSU0_ERR_CTRL_FLD_RESERVED_1_WIDTH 9
`define DDRMC5_NOC_NSU0_ERR_CTRL_WIDTH 23

/* NSU1_ERR_CTRL */
`define DDRMC5_NOC_NSU1_ERR_CTRL_OFFSET 17'h5f4
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_RESERVED 11:0
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_PAR_RESP_ERR_EN 12
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_PAR_RESP_ERR_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_FATAL_DROP_EN 13
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_FATAL_DROP_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_SEL 15:14
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_SEL_WIDTH 2
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_DW_EN 16
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_DW_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_CW_EN 17
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_CW_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_R_EN 18
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_R_EN_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_DW_DONE 19
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_DW_DONE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_CW_DONE 20
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_CW_DONE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_R_DONE 21
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_R_DONE_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_PERSISTENT 22
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_PERSISTENT_WIDTH 1
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_RESERVED_1 31:23
`define DDRMC5_NOC_NSU1_ERR_CTRL_FLD_RESERVED_1_WIDTH 9
`define DDRMC5_NOC_NSU1_ERR_CTRL_WIDTH 23

/* ECC_ERR_INJ_NSU0 */
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_OFFSET 17'h5f8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_BIT_0 7:0
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_BIT_0_WIDTH 8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_BIT_1 15:8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_BIT_1_WIDTH 8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_EN_RD 16
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_EN_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_DONE_RD 17
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_DONE_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_EN_WR 18
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_EN_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_DONE_WR 19
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_ECC_DONE_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_EN_RD 20
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_EN_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_DONE_RD 21
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_DONE_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_EN_WR 22
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_EN_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_DONE_WR 23
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_DST_PAR_DONE_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_PERSISTENT 24
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_PERSISTENT_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_RESERVED 31:25
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_ECC_ERR_INJ_NSU0_WIDTH 25

/* ECC_ERR_INJ_NSU1 */
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_OFFSET 17'h5fc
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_BIT_0 7:0
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_BIT_0_WIDTH 8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_BIT_1 15:8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_BIT_1_WIDTH 8
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_EN_RD 16
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_EN_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_DONE_RD 17
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_DONE_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_EN_WR 18
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_EN_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_DONE_WR 19
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_ECC_DONE_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_EN_RD 20
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_EN_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_DONE_RD 21
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_DONE_RD_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_EN_WR 22
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_EN_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_DONE_WR 23
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_DST_PAR_DONE_WR_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_PERSISTENT 24
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_PERSISTENT_WIDTH 1
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_RESERVED 31:25
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_FLD_RESERVED_WIDTH 7
`define DDRMC5_NOC_ECC_ERR_INJ_NSU1_WIDTH 25

/* ILA_MUX_P0_N0 */
`define DDRMC5_NOC_ILA_MUX_P0_N0_OFFSET 17'h600
`define DDRMC5_NOC_ILA_MUX_P0_N0_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N0_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N0_WIDTH 32

/* ILA_MUX_P0_N1 */
`define DDRMC5_NOC_ILA_MUX_P0_N1_OFFSET 17'h604
`define DDRMC5_NOC_ILA_MUX_P0_N1_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N1_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N1_WIDTH 32

/* ILA_MUX_P0_N2 */
`define DDRMC5_NOC_ILA_MUX_P0_N2_OFFSET 17'h608
`define DDRMC5_NOC_ILA_MUX_P0_N2_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N2_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N2_WIDTH 32

/* ILA_MUX_P0_N3 */
`define DDRMC5_NOC_ILA_MUX_P0_N3_OFFSET 17'h60c
`define DDRMC5_NOC_ILA_MUX_P0_N3_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N3_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N3_WIDTH 32

/* ILA_MUX_P0_N4 */
`define DDRMC5_NOC_ILA_MUX_P0_N4_OFFSET 17'h610
`define DDRMC5_NOC_ILA_MUX_P0_N4_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N4_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N4_WIDTH 32

/* ILA_MUX_P0_N5 */
`define DDRMC5_NOC_ILA_MUX_P0_N5_OFFSET 17'h614
`define DDRMC5_NOC_ILA_MUX_P0_N5_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N5_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N5_WIDTH 32

/* ILA_MUX_P0_N6 */
`define DDRMC5_NOC_ILA_MUX_P0_N6_OFFSET 17'h618
`define DDRMC5_NOC_ILA_MUX_P0_N6_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N6_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N6_WIDTH 32

/* ILA_MUX_P0_N7 */
`define DDRMC5_NOC_ILA_MUX_P0_N7_OFFSET 17'h61c
`define DDRMC5_NOC_ILA_MUX_P0_N7_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N7_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N7_WIDTH 32

/* ILA_MUX_P0_N8 */
`define DDRMC5_NOC_ILA_MUX_P0_N8_OFFSET 17'h620
`define DDRMC5_NOC_ILA_MUX_P0_N8_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N8_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N8_WIDTH 32

/* ILA_MUX_P0_N9 */
`define DDRMC5_NOC_ILA_MUX_P0_N9_OFFSET 17'h624
`define DDRMC5_NOC_ILA_MUX_P0_N9_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N9_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N9_WIDTH 32

/* ILA_MUX_P0_N10 */
`define DDRMC5_NOC_ILA_MUX_P0_N10_OFFSET 17'h628
`define DDRMC5_NOC_ILA_MUX_P0_N10_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N10_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N10_WIDTH 32

/* ILA_MUX_P0_N11 */
`define DDRMC5_NOC_ILA_MUX_P0_N11_OFFSET 17'h62c
`define DDRMC5_NOC_ILA_MUX_P0_N11_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N11_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N11_WIDTH 32

/* ILA_MUX_P0_N12 */
`define DDRMC5_NOC_ILA_MUX_P0_N12_OFFSET 17'h630
`define DDRMC5_NOC_ILA_MUX_P0_N12_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N12_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N12_WIDTH 32

/* ILA_MUX_P0_N13 */
`define DDRMC5_NOC_ILA_MUX_P0_N13_OFFSET 17'h634
`define DDRMC5_NOC_ILA_MUX_P0_N13_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N13_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N13_WIDTH 32

/* ILA_MUX_P0_N14 */
`define DDRMC5_NOC_ILA_MUX_P0_N14_OFFSET 17'h638
`define DDRMC5_NOC_ILA_MUX_P0_N14_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N14_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N14_WIDTH 32

/* ILA_MUX_P0_N15 */
`define DDRMC5_NOC_ILA_MUX_P0_N15_OFFSET 17'h63c
`define DDRMC5_NOC_ILA_MUX_P0_N15_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N15_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N15_WIDTH 32

/* ILA_MUX_P0_N16 */
`define DDRMC5_NOC_ILA_MUX_P0_N16_OFFSET 17'h640
`define DDRMC5_NOC_ILA_MUX_P0_N16_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N16_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N16_WIDTH 32

/* ILA_MUX_P0_N17 */
`define DDRMC5_NOC_ILA_MUX_P0_N17_OFFSET 17'h644
`define DDRMC5_NOC_ILA_MUX_P0_N17_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N17_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N17_WIDTH 32

/* ILA_MUX_P0_N18 */
`define DDRMC5_NOC_ILA_MUX_P0_N18_OFFSET 17'h648
`define DDRMC5_NOC_ILA_MUX_P0_N18_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N18_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N18_WIDTH 32

/* ILA_MUX_P0_N19 */
`define DDRMC5_NOC_ILA_MUX_P0_N19_OFFSET 17'h64c
`define DDRMC5_NOC_ILA_MUX_P0_N19_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N19_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N19_WIDTH 32

/* ILA_MUX_P0_N20 */
`define DDRMC5_NOC_ILA_MUX_P0_N20_OFFSET 17'h650
`define DDRMC5_NOC_ILA_MUX_P0_N20_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P0_N20_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P0_N20_WIDTH 32

/* ILA_MUX_P1_N0 */
`define DDRMC5_NOC_ILA_MUX_P1_N0_OFFSET 17'h654
`define DDRMC5_NOC_ILA_MUX_P1_N0_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N0_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N0_WIDTH 32

/* ILA_MUX_P1_N1 */
`define DDRMC5_NOC_ILA_MUX_P1_N1_OFFSET 17'h658
`define DDRMC5_NOC_ILA_MUX_P1_N1_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N1_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N1_WIDTH 32

/* ILA_MUX_P1_N2 */
`define DDRMC5_NOC_ILA_MUX_P1_N2_OFFSET 17'h65c
`define DDRMC5_NOC_ILA_MUX_P1_N2_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N2_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N2_WIDTH 32

/* ILA_MUX_P1_N3 */
`define DDRMC5_NOC_ILA_MUX_P1_N3_OFFSET 17'h660
`define DDRMC5_NOC_ILA_MUX_P1_N3_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N3_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N3_WIDTH 32

/* ILA_MUX_P1_N4 */
`define DDRMC5_NOC_ILA_MUX_P1_N4_OFFSET 17'h664
`define DDRMC5_NOC_ILA_MUX_P1_N4_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N4_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N4_WIDTH 32

/* ILA_MUX_P1_N5 */
`define DDRMC5_NOC_ILA_MUX_P1_N5_OFFSET 17'h668
`define DDRMC5_NOC_ILA_MUX_P1_N5_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N5_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N5_WIDTH 32

/* ILA_MUX_P1_N6 */
`define DDRMC5_NOC_ILA_MUX_P1_N6_OFFSET 17'h66c
`define DDRMC5_NOC_ILA_MUX_P1_N6_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N6_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N6_WIDTH 32

/* ILA_MUX_P1_N7 */
`define DDRMC5_NOC_ILA_MUX_P1_N7_OFFSET 17'h670
`define DDRMC5_NOC_ILA_MUX_P1_N7_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N7_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N7_WIDTH 32

/* ILA_MUX_P1_N8 */
`define DDRMC5_NOC_ILA_MUX_P1_N8_OFFSET 17'h674
`define DDRMC5_NOC_ILA_MUX_P1_N8_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N8_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N8_WIDTH 32

/* ILA_MUX_P1_N9 */
`define DDRMC5_NOC_ILA_MUX_P1_N9_OFFSET 17'h678
`define DDRMC5_NOC_ILA_MUX_P1_N9_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N9_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N9_WIDTH 32

/* ILA_MUX_P1_N10 */
`define DDRMC5_NOC_ILA_MUX_P1_N10_OFFSET 17'h67c
`define DDRMC5_NOC_ILA_MUX_P1_N10_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N10_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N10_WIDTH 32

/* ILA_MUX_P1_N11 */
`define DDRMC5_NOC_ILA_MUX_P1_N11_OFFSET 17'h680
`define DDRMC5_NOC_ILA_MUX_P1_N11_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N11_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N11_WIDTH 32

/* ILA_MUX_P1_N12 */
`define DDRMC5_NOC_ILA_MUX_P1_N12_OFFSET 17'h684
`define DDRMC5_NOC_ILA_MUX_P1_N12_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N12_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N12_WIDTH 32

/* ILA_MUX_P1_N13 */
`define DDRMC5_NOC_ILA_MUX_P1_N13_OFFSET 17'h688
`define DDRMC5_NOC_ILA_MUX_P1_N13_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N13_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N13_WIDTH 32

/* ILA_MUX_P1_N14 */
`define DDRMC5_NOC_ILA_MUX_P1_N14_OFFSET 17'h68c
`define DDRMC5_NOC_ILA_MUX_P1_N14_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N14_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N14_WIDTH 32

/* ILA_MUX_P1_N15 */
`define DDRMC5_NOC_ILA_MUX_P1_N15_OFFSET 17'h690
`define DDRMC5_NOC_ILA_MUX_P1_N15_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N15_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N15_WIDTH 32

/* ILA_MUX_P1_N16 */
`define DDRMC5_NOC_ILA_MUX_P1_N16_OFFSET 17'h694
`define DDRMC5_NOC_ILA_MUX_P1_N16_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N16_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N16_WIDTH 32

/* ILA_MUX_P1_N17 */
`define DDRMC5_NOC_ILA_MUX_P1_N17_OFFSET 17'h698
`define DDRMC5_NOC_ILA_MUX_P1_N17_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N17_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N17_WIDTH 32

/* ILA_MUX_P1_N18 */
`define DDRMC5_NOC_ILA_MUX_P1_N18_OFFSET 17'h69c
`define DDRMC5_NOC_ILA_MUX_P1_N18_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N18_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N18_WIDTH 32

/* ILA_MUX_P1_N19 */
`define DDRMC5_NOC_ILA_MUX_P1_N19_OFFSET 17'h6a0
`define DDRMC5_NOC_ILA_MUX_P1_N19_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N19_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N19_WIDTH 32

/* ILA_MUX_P1_N20 */
`define DDRMC5_NOC_ILA_MUX_P1_N20_OFFSET 17'h6a4
`define DDRMC5_NOC_ILA_MUX_P1_N20_FLD_DBG_MC_SEL 31:0
`define DDRMC5_NOC_ILA_MUX_P1_N20_FLD_DBG_MC_SEL_WIDTH 32
`define DDRMC5_NOC_ILA_MUX_P1_N20_WIDTH 32

/* NA_ERR_CTRL_0 */
`define DDRMC5_NOC_NA_ERR_CTRL_0_OFFSET 17'h6a8
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_RESERVED 27:0
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_DROP_PAR_ERR_EN 28
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_DROP_PAR_ERR_EN_WIDTH 1
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_RESERVED_1 31:29
`define DDRMC5_NOC_NA_ERR_CTRL_0_FLD_RESERVED_1_WIDTH 3
`define DDRMC5_NOC_NA_ERR_CTRL_0_WIDTH 29

/* REG_DBG_MUX_SEL */
`define DDRMC5_NOC_REG_DBG_MUX_SEL_OFFSET 17'h6ac
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_OUT_SEL 0
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_OUT_SEL_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_IN_SEL 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_IN_SEL_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_DBG_EN 2
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_DBG_EN_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_TRIG_EN 3
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_TRIG_EN_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_CLK_DIV 4
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_CLK_DIV_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_POST_TRIG_CNT 7:5
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_POST_TRIG_CNT_WIDTH 3
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_DAT_DISC 8
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_DAT_DISC_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_TRIG_DONE 9
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_TRIG_DONE_WIDTH 1
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_RESERVED 31:10
`define DDRMC5_NOC_REG_DBG_MUX_SEL_FLD_RESERVED_WIDTH 22
`define DDRMC5_NOC_REG_DBG_MUX_SEL_WIDTH 10

/* REG_DBG_DATA_SEL */
`define DDRMC5_NOC_REG_DBG_DATA_SEL_OFFSET 17'h6b0
`define DDRMC5_NOC_REG_DBG_DATA_SEL_FLD_DDRMC 7:0
`define DDRMC5_NOC_REG_DBG_DATA_SEL_FLD_DDRMC_WIDTH 8
`define DDRMC5_NOC_REG_DBG_DATA_SEL_FLD_RESERVED 31:8
`define DDRMC5_NOC_REG_DBG_DATA_SEL_FLD_RESERVED_WIDTH 24
`define DDRMC5_NOC_REG_DBG_DATA_SEL_WIDTH 8

/* REG_DBG_TRIG_MVAL_L */
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_L_OFFSET 17'h6b4
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_L_FLD_DDRMC 31:0
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_L_FLD_DDRMC_WIDTH 32
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_L_WIDTH 32

/* REG_DBG_TRIG_MVAL_U */
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_U_OFFSET 17'h6b8
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_U_FLD_DDRMC 31:0
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_U_FLD_DDRMC_WIDTH 32
`define DDRMC5_NOC_REG_DBG_TRIG_MVAL_U_WIDTH 32

/* REG_DBG_TRIG_MASK_L */
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_L_OFFSET 17'h6bc
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_L_FLD_DDRMC 31:0
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_L_FLD_DDRMC_WIDTH 32
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_L_WIDTH 32

/* REG_DBG_TRIG_MASK_U */
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_U_OFFSET 17'h6c0
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_U_FLD_DDRMC 31:0
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_U_FLD_DDRMC_WIDTH 32
`define DDRMC5_NOC_REG_DBG_TRIG_MASK_U_WIDTH 32

/* DDRMC_CLK_MUX */
`define DDRMC5_NOC_DDRMC_CLK_MUX_OFFSET 17'h6c4
`define DDRMC5_NOC_DDRMC_CLK_MUX_FLD_SEL 0
`define DDRMC5_NOC_DDRMC_CLK_MUX_FLD_SEL_WIDTH 1
`define DDRMC5_NOC_DDRMC_CLK_MUX_FLD_RESERVED 31:1
`define DDRMC5_NOC_DDRMC_CLK_MUX_FLD_RESERVED_WIDTH 31
`define DDRMC5_NOC_DDRMC_CLK_MUX_WIDTH 1

/* XMPU_CRPTO_CFG0_0 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_OFFSET 17'h10000
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_0_WIDTH 8

/* XMPU_CRPTO_CFG1_0 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_OFFSET 17'h10004
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_0_WIDTH 28

/* XMPU_CRPTO_CFG2_0 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_OFFSET 17'h10008
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_0_WIDTH 28

/* XMPU_CRPTO_CFG0_1 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_OFFSET 17'h1000c
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_1_WIDTH 8

/* XMPU_CRPTO_CFG1_1 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_OFFSET 17'h10010
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_1_WIDTH 28

/* XMPU_CRPTO_CFG2_1 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_OFFSET 17'h10014
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_1_WIDTH 28

/* XMPU_CRPTO_CFG0_2 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_OFFSET 17'h10018
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_2_WIDTH 8

/* XMPU_CRPTO_CFG1_2 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_OFFSET 17'h1001c
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_2_WIDTH 28

/* XMPU_CRPTO_CFG2_2 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_OFFSET 17'h10020
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_2_WIDTH 28

/* XMPU_CRPTO_CFG0_3 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_OFFSET 17'h10024
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_3_WIDTH 8

/* XMPU_CRPTO_CFG1_3 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_OFFSET 17'h10028
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_3_WIDTH 28

/* XMPU_CRPTO_CFG2_3 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_OFFSET 17'h1002c
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_3_WIDTH 28

/* XMPU_CRPTO_CFG0_4 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_OFFSET 17'h10030
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_4_WIDTH 8

/* XMPU_CRPTO_CFG1_4 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_OFFSET 17'h10034
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_4_WIDTH 28

/* XMPU_CRPTO_CFG2_4 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_OFFSET 17'h10038
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_4_WIDTH 28

/* XMPU_CRPTO_CFG0_5 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_OFFSET 17'h1003c
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_5_WIDTH 8

/* XMPU_CRPTO_CFG1_5 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_OFFSET 17'h10040
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_5_WIDTH 28

/* XMPU_CRPTO_CFG2_5 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_OFFSET 17'h10044
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_5_WIDTH 28

/* XMPU_CRPTO_CFG0_6 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_OFFSET 17'h10048
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_6_WIDTH 8

/* XMPU_CRPTO_CFG1_6 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_OFFSET 17'h1004c
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_6_WIDTH 28

/* XMPU_CRPTO_CFG2_6 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_OFFSET 17'h10050
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_6_WIDTH 28

/* XMPU_CRPTO_CFG0_7 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_OFFSET 17'h10054
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_7_WIDTH 8

/* XMPU_CRPTO_CFG1_7 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_OFFSET 17'h10058
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_7_WIDTH 28

/* XMPU_CRPTO_CFG2_7 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_OFFSET 17'h1005c
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_7_WIDTH 28

/* XMPU_CRPTO_CFG0_8 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_OFFSET 17'h10060
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_8_WIDTH 8

/* XMPU_CRPTO_CFG1_8 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_OFFSET 17'h10064
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_8_WIDTH 28

/* XMPU_CRPTO_CFG2_8 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_OFFSET 17'h10068
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_8_WIDTH 28

/* XMPU_CRPTO_CFG0_9 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_OFFSET 17'h1006c
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_9_WIDTH 8

/* XMPU_CRPTO_CFG1_9 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_OFFSET 17'h10070
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_9_WIDTH 28

/* XMPU_CRPTO_CFG2_9 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_OFFSET 17'h10074
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_9_WIDTH 28

/* XMPU_CRPTO_CFG0_10 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_OFFSET 17'h10078
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_10_WIDTH 8

/* XMPU_CRPTO_CFG1_10 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_OFFSET 17'h1007c
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_10_WIDTH 28

/* XMPU_CRPTO_CFG2_10 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_OFFSET 17'h10080
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_10_WIDTH 28

/* XMPU_CRPTO_CFG0_11 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_OFFSET 17'h10084
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_11_WIDTH 8

/* XMPU_CRPTO_CFG1_11 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_OFFSET 17'h10088
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_11_WIDTH 28

/* XMPU_CRPTO_CFG2_11 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_OFFSET 17'h1008c
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_11_WIDTH 28

/* XMPU_CRPTO_CFG0_12 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_OFFSET 17'h10090
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_12_WIDTH 8

/* XMPU_CRPTO_CFG1_12 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_OFFSET 17'h10094
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_12_WIDTH 28

/* XMPU_CRPTO_CFG2_12 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_OFFSET 17'h10098
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_12_WIDTH 28

/* XMPU_CRPTO_CFG0_13 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_OFFSET 17'h1009c
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_13_WIDTH 8

/* XMPU_CRPTO_CFG1_13 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_OFFSET 17'h100a0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_13_WIDTH 28

/* XMPU_CRPTO_CFG2_13 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_OFFSET 17'h100a4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_13_WIDTH 28

/* XMPU_CRPTO_CFG0_14 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_OFFSET 17'h100a8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_14_WIDTH 8

/* XMPU_CRPTO_CFG1_14 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_OFFSET 17'h100ac
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_14_WIDTH 28

/* XMPU_CRPTO_CFG2_14 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_OFFSET 17'h100b0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_14_WIDTH 28

/* XMPU_CRPTO_CFG0_15 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_OFFSET 17'h100b4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_ENC_TYPE 1:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_ENC_TYPE_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_RESERVED 3:2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_NUM_KEY 7:4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_NUM_KEY_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_RESERVED_1 31:8
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_FLD_RESERVED_1_WIDTH 24
`define DDRMC5_NOC_XMPU_CRPTO_CFG0_15_WIDTH 8

/* XMPU_CRPTO_CFG1_15 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_OFFSET 17'h100b8
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_FLD_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_FLD_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG1_15_WIDTH 28

/* XMPU_CRPTO_CFG2_15 */
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_OFFSET 17'h100bc
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_FLD_ABS_MAX_KEY_USAGE 27:0
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_FLD_ABS_MAX_KEY_USAGE_WIDTH 28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_FLD_RESERVED 31:28
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_XMPU_CRPTO_CFG2_15_WIDTH 28

/* REG_ADEC0 */
`define DDRMC5_NOC_REG_ADEC0_OFFSET 17'h100c0
`define DDRMC5_NOC_REG_ADEC0_FLD_LOW_MEM_BASE 19:0
`define DDRMC5_NOC_REG_ADEC0_FLD_LOW_MEM_BASE_WIDTH 20
`define DDRMC5_NOC_REG_ADEC0_FLD_RESERVED 31:20
`define DDRMC5_NOC_REG_ADEC0_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_REG_ADEC0_WIDTH 20

/* REG_ADEC1 */
`define DDRMC5_NOC_REG_ADEC1_OFFSET 17'h100c4
`define DDRMC5_NOC_REG_ADEC1_FLD_LOW_MEM_OFFSET 19:0
`define DDRMC5_NOC_REG_ADEC1_FLD_LOW_MEM_OFFSET_WIDTH 20
`define DDRMC5_NOC_REG_ADEC1_FLD_RESERVED 31:20
`define DDRMC5_NOC_REG_ADEC1_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_REG_ADEC1_WIDTH 20

/* REG_ADEC2 */
`define DDRMC5_NOC_REG_ADEC2_OFFSET 17'h100c8
`define DDRMC5_NOC_REG_ADEC2_FLD_HIGH_MEM_BASE 19:0
`define DDRMC5_NOC_REG_ADEC2_FLD_HIGH_MEM_BASE_WIDTH 20
`define DDRMC5_NOC_REG_ADEC2_FLD_HIGH_MEM_EN 20
`define DDRMC5_NOC_REG_ADEC2_FLD_HIGH_MEM_EN_WIDTH 1
`define DDRMC5_NOC_REG_ADEC2_FLD_RESERVED 31:21
`define DDRMC5_NOC_REG_ADEC2_FLD_RESERVED_WIDTH 11
`define DDRMC5_NOC_REG_ADEC2_WIDTH 21

/* REG_ADEC3 */
`define DDRMC5_NOC_REG_ADEC3_OFFSET 17'h100cc
`define DDRMC5_NOC_REG_ADEC3_FLD_HIGH_MEM_OFFSET 19:0
`define DDRMC5_NOC_REG_ADEC3_FLD_HIGH_MEM_OFFSET_WIDTH 20
`define DDRMC5_NOC_REG_ADEC3_FLD_RESERVED 31:20
`define DDRMC5_NOC_REG_ADEC3_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_REG_ADEC3_WIDTH 20

/* REG_ADEC4 */
`define DDRMC5_NOC_REG_ADEC4_OFFSET 17'h100d0
`define DDRMC5_NOC_REG_ADEC4_FLD_RANK_0 5:0
`define DDRMC5_NOC_REG_ADEC4_FLD_RANK_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC4_FLD_RANK_1 11:6
`define DDRMC5_NOC_REG_ADEC4_FLD_RANK_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC4_FLD_RESERVED 31:12
`define DDRMC5_NOC_REG_ADEC4_FLD_RESERVED_WIDTH 20
`define DDRMC5_NOC_REG_ADEC4_WIDTH 12

/* REG_ADEC5 */
`define DDRMC5_NOC_REG_ADEC5_OFFSET 17'h100d4
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_0 5:0
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_1 11:6
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_2 17:12
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_2_WIDTH 6
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_3 23:18
`define DDRMC5_NOC_REG_ADEC5_FLD_LRANK_3_WIDTH 6
`define DDRMC5_NOC_REG_ADEC5_FLD_RESERVED 31:24
`define DDRMC5_NOC_REG_ADEC5_FLD_RESERVED_WIDTH 8
`define DDRMC5_NOC_REG_ADEC5_WIDTH 24

/* REG_ADEC6 */
`define DDRMC5_NOC_REG_ADEC6_OFFSET 17'h100d8
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_0 5:0
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_1 11:6
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_2 17:12
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_2_WIDTH 6
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_3 23:18
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_3_WIDTH 6
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_4 29:24
`define DDRMC5_NOC_REG_ADEC6_FLD_ROW_4_WIDTH 6
`define DDRMC5_NOC_REG_ADEC6_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC6_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC6_WIDTH 30

/* REG_ADEC7 */
`define DDRMC5_NOC_REG_ADEC7_OFFSET 17'h100dc
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_5 5:0
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_5_WIDTH 6
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_6 11:6
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_6_WIDTH 6
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_7 17:12
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_7_WIDTH 6
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_8 23:18
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_8_WIDTH 6
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_9 29:24
`define DDRMC5_NOC_REG_ADEC7_FLD_ROW_9_WIDTH 6
`define DDRMC5_NOC_REG_ADEC7_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC7_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC7_WIDTH 30

/* REG_ADEC8 */
`define DDRMC5_NOC_REG_ADEC8_OFFSET 17'h100e0
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_10 5:0
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_10_WIDTH 6
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_11 11:6
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_11_WIDTH 6
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_12 17:12
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_12_WIDTH 6
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_13 23:18
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_13_WIDTH 6
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_14 29:24
`define DDRMC5_NOC_REG_ADEC8_FLD_ROW_14_WIDTH 6
`define DDRMC5_NOC_REG_ADEC8_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC8_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC8_WIDTH 30

/* REG_ADEC9 */
`define DDRMC5_NOC_REG_ADEC9_OFFSET 17'h100e4
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_15 5:0
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_15_WIDTH 6
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_16 11:6
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_16_WIDTH 6
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_17 17:12
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_17_WIDTH 6
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_18 23:18
`define DDRMC5_NOC_REG_ADEC9_FLD_ROW_18_WIDTH 6
`define DDRMC5_NOC_REG_ADEC9_FLD_COL_0 29:24
`define DDRMC5_NOC_REG_ADEC9_FLD_COL_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC9_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC9_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC9_WIDTH 30

/* REG_ADEC10 */
`define DDRMC5_NOC_REG_ADEC10_OFFSET 17'h100e8
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_1 5:0
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_2 11:6
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_2_WIDTH 6
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_3 17:12
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_3_WIDTH 6
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_4 23:18
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_4_WIDTH 6
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_5 29:24
`define DDRMC5_NOC_REG_ADEC10_FLD_COL_5_WIDTH 6
`define DDRMC5_NOC_REG_ADEC10_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC10_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC10_WIDTH 30

/* REG_ADEC11 */
`define DDRMC5_NOC_REG_ADEC11_OFFSET 17'h100ec
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_6 5:0
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_6_WIDTH 6
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_7 11:6
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_7_WIDTH 6
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_8 17:12
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_8_WIDTH 6
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_9 23:18
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_9_WIDTH 6
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_10 29:24
`define DDRMC5_NOC_REG_ADEC11_FLD_COL_10_WIDTH 6
`define DDRMC5_NOC_REG_ADEC11_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC11_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC11_WIDTH 30

/* REG_ADEC12 */
`define DDRMC5_NOC_REG_ADEC12_OFFSET 17'h100f0
`define DDRMC5_NOC_REG_ADEC12_FLD_BANK_0 5:0
`define DDRMC5_NOC_REG_ADEC12_FLD_BANK_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC12_FLD_BANK_1 11:6
`define DDRMC5_NOC_REG_ADEC12_FLD_BANK_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_0 17:12
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_1 23:18
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_2 29:24
`define DDRMC5_NOC_REG_ADEC12_FLD_GROUP_2_WIDTH 6
`define DDRMC5_NOC_REG_ADEC12_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC12_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC12_WIDTH 30

/* REG_ADEC13 */
`define DDRMC5_NOC_REG_ADEC13_OFFSET 17'h100f4
`define DDRMC5_NOC_REG_ADEC13_FLD_INTERLEAVE_SEL 3:0
`define DDRMC5_NOC_REG_ADEC13_FLD_INTERLEAVE_SEL_WIDTH 4
`define DDRMC5_NOC_REG_ADEC13_FLD_INTERLEAVE_SIZE 6:4
`define DDRMC5_NOC_REG_ADEC13_FLD_INTERLEAVE_SIZE_WIDTH 3
`define DDRMC5_NOC_REG_ADEC13_FLD_RESERVED 31:7
`define DDRMC5_NOC_REG_ADEC13_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_REG_ADEC13_WIDTH 7

/* REG_ADEC14 */
`define DDRMC5_NOC_REG_ADEC14_OFFSET 17'h100f8
`define DDRMC5_NOC_REG_ADEC14_FLD_ILC_MEM_BASE 27:0
`define DDRMC5_NOC_REG_ADEC14_FLD_ILC_MEM_BASE_WIDTH 28
`define DDRMC5_NOC_REG_ADEC14_FLD_ILC_HIGN_MEM_EN 28
`define DDRMC5_NOC_REG_ADEC14_FLD_ILC_HIGN_MEM_EN_WIDTH 1
`define DDRMC5_NOC_REG_ADEC14_FLD_RESERVED 31:29
`define DDRMC5_NOC_REG_ADEC14_FLD_RESERVED_WIDTH 3
`define DDRMC5_NOC_REG_ADEC14_WIDTH 29

/* REG_ADEC15 */
`define DDRMC5_NOC_REG_ADEC15_OFFSET 17'h100fc
`define DDRMC5_NOC_REG_ADEC15_FLD_ILC_MEM_SIZE 27:0
`define DDRMC5_NOC_REG_ADEC15_FLD_ILC_MEM_SIZE_WIDTH 28
`define DDRMC5_NOC_REG_ADEC15_FLD_RESERVED 31:28
`define DDRMC5_NOC_REG_ADEC15_FLD_RESERVED_WIDTH 4
`define DDRMC5_NOC_REG_ADEC15_WIDTH 28

/* REG_ADEC16 */
`define DDRMC5_NOC_REG_ADEC16_OFFSET 17'h10100
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_ECC_STORAGE_BASE 27:0
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_ECC_STORAGE_BASE_WIDTH 28
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_ECC_HIGN_EN 28
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_ECC_HIGN_EN_WIDTH 1
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_BYPASS_EN 29
`define DDRMC5_NOC_REG_ADEC16_FLD_ILC_BYPASS_EN_WIDTH 1
`define DDRMC5_NOC_REG_ADEC16_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC16_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC16_WIDTH 30

/* REG_ADEC_ILC */
`define DDRMC5_NOC_REG_ADEC_ILC_OFFSET 17'h10104
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_0 5:0
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_0_WIDTH 6
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_1 11:6
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_1_WIDTH 6
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_2 17:12
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_ECC_COL_2_WIDTH 6
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_RESERVED 31:30
`define DDRMC5_NOC_REG_ADEC_ILC_FLD_RESERVED_WIDTH 2
`define DDRMC5_NOC_REG_ADEC_ILC_WIDTH 18

/* REG_ADEC_MEMFILL0_LOW */
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_LOW_OFFSET 17'h10108
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_LOW_FLD_BASE 31:0
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_LOW_FLD_BASE_WIDTH 32
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_LOW_WIDTH 32

/* REG_ADEC_MEMFILL1_LOW */
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_LOW_OFFSET 17'h1010c
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_LOW_FLD_RANGE 31:0
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_LOW_FLD_RANGE_WIDTH 32
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_LOW_WIDTH 32

/* REG_ADEC_MEMFILL0_HIGH */
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_HIGH_OFFSET 17'h10110
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_HIGH_FLD_BASE 31:0
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_HIGH_FLD_BASE_WIDTH 32
`define DDRMC5_NOC_REG_ADEC_MEMFILL0_HIGH_WIDTH 32

/* REG_ADEC_MEMFILL1_HIGH */
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_HIGH_OFFSET 17'h10114
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_HIGH_FLD_RANGE 31:0
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_HIGH_FLD_RANGE_WIDTH 32
`define DDRMC5_NOC_REG_ADEC_MEMFILL1_HIGH_WIDTH 32

/* XMPU_CTRL */
`define DDRMC5_NOC_XMPU_CTRL_OFFSET 17'h12000
`define DDRMC5_NOC_XMPU_CTRL_FLD_DEFRDALLOWED 0
`define DDRMC5_NOC_XMPU_CTRL_FLD_DEFRDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_DEFWRALLOWED 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_DEFWRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_HIDEALLOWED 2
`define DDRMC5_NOC_XMPU_CTRL_FLD_HIDEALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_ALIGNCFG 3
`define DDRMC5_NOC_XMPU_CTRL_FLD_ALIGNCFG_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_RDPERMVIO_MASK 4
`define DDRMC5_NOC_XMPU_CTRL_FLD_RDPERMVIO_MASK_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_WRPERMVIO_MASK 5
`define DDRMC5_NOC_XMPU_CTRL_FLD_WRPERMVIO_MASK_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_SECURITYVIO_MASK 6
`define DDRMC5_NOC_XMPU_CTRL_FLD_SECURITYVIO_MASK_WIDTH 1
`define DDRMC5_NOC_XMPU_CTRL_FLD_RESERVED 31:7
`define DDRMC5_NOC_XMPU_CTRL_FLD_RESERVED_WIDTH 25
`define DDRMC5_NOC_XMPU_CTRL_WIDTH 7

/* XMPU_START_LO0 */
`define DDRMC5_NOC_XMPU_START_LO0_OFFSET 17'h12004
`define DDRMC5_NOC_XMPU_START_LO0_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO0_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO0_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO0_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO0_WIDTH 32

/* XMPU_START_HI0 */
`define DDRMC5_NOC_XMPU_START_HI0_OFFSET 17'h12008
`define DDRMC5_NOC_XMPU_START_HI0_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI0_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI0_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI0_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI0_WIDTH 16

/* XMPU_END_LO0 */
`define DDRMC5_NOC_XMPU_END_LO0_OFFSET 17'h1200c
`define DDRMC5_NOC_XMPU_END_LO0_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO0_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO0_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO0_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO0_WIDTH 32

/* XMPU_END_HI0 */
`define DDRMC5_NOC_XMPU_END_HI0_OFFSET 17'h12010
`define DDRMC5_NOC_XMPU_END_HI0_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI0_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI0_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI0_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI0_WIDTH 16

/* XMPU_MASTER0 */
`define DDRMC5_NOC_XMPU_MASTER0_OFFSET 17'h12014
`define DDRMC5_NOC_XMPU_MASTER0_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER0_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER0_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER0_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER0_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER0_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER0_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER0_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER0_WIDTH 26

/* XMPU_CONFIG0 */
`define DDRMC5_NOC_XMPU_CONFIG0_OFFSET 17'h12018
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG0_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG0_WIDTH 5

/* XMPU_START_LO1 */
`define DDRMC5_NOC_XMPU_START_LO1_OFFSET 17'h1201c
`define DDRMC5_NOC_XMPU_START_LO1_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO1_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO1_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO1_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO1_WIDTH 32

/* XMPU_START_HI1 */
`define DDRMC5_NOC_XMPU_START_HI1_OFFSET 17'h12020
`define DDRMC5_NOC_XMPU_START_HI1_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI1_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI1_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI1_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI1_WIDTH 16

/* XMPU_END_LO1 */
`define DDRMC5_NOC_XMPU_END_LO1_OFFSET 17'h12024
`define DDRMC5_NOC_XMPU_END_LO1_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO1_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO1_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO1_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO1_WIDTH 32

/* XMPU_END_HI1 */
`define DDRMC5_NOC_XMPU_END_HI1_OFFSET 17'h12028
`define DDRMC5_NOC_XMPU_END_HI1_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI1_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI1_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI1_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI1_WIDTH 16

/* XMPU_MASTER1 */
`define DDRMC5_NOC_XMPU_MASTER1_OFFSET 17'h1202c
`define DDRMC5_NOC_XMPU_MASTER1_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER1_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER1_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER1_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER1_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER1_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER1_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER1_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER1_WIDTH 26

/* XMPU_CONFIG1 */
`define DDRMC5_NOC_XMPU_CONFIG1_OFFSET 17'h12030
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG1_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG1_WIDTH 5

/* XMPU_START_LO2 */
`define DDRMC5_NOC_XMPU_START_LO2_OFFSET 17'h12034
`define DDRMC5_NOC_XMPU_START_LO2_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO2_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO2_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO2_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO2_WIDTH 32

/* XMPU_START_HI2 */
`define DDRMC5_NOC_XMPU_START_HI2_OFFSET 17'h12038
`define DDRMC5_NOC_XMPU_START_HI2_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI2_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI2_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI2_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI2_WIDTH 16

/* XMPU_END_LO2 */
`define DDRMC5_NOC_XMPU_END_LO2_OFFSET 17'h1203c
`define DDRMC5_NOC_XMPU_END_LO2_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO2_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO2_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO2_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO2_WIDTH 32

/* XMPU_END_HI2 */
`define DDRMC5_NOC_XMPU_END_HI2_OFFSET 17'h12040
`define DDRMC5_NOC_XMPU_END_HI2_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI2_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI2_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI2_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI2_WIDTH 16

/* XMPU_MASTER2 */
`define DDRMC5_NOC_XMPU_MASTER2_OFFSET 17'h12044
`define DDRMC5_NOC_XMPU_MASTER2_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER2_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER2_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER2_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER2_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER2_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER2_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER2_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER2_WIDTH 26

/* XMPU_CONFIG2 */
`define DDRMC5_NOC_XMPU_CONFIG2_OFFSET 17'h12048
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG2_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG2_WIDTH 5

/* XMPU_START_LO3 */
`define DDRMC5_NOC_XMPU_START_LO3_OFFSET 17'h1204c
`define DDRMC5_NOC_XMPU_START_LO3_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO3_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO3_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO3_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO3_WIDTH 32

/* XMPU_START_HI3 */
`define DDRMC5_NOC_XMPU_START_HI3_OFFSET 17'h12050
`define DDRMC5_NOC_XMPU_START_HI3_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI3_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI3_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI3_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI3_WIDTH 16

/* XMPU_END_LO3 */
`define DDRMC5_NOC_XMPU_END_LO3_OFFSET 17'h12054
`define DDRMC5_NOC_XMPU_END_LO3_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO3_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO3_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO3_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO3_WIDTH 32

/* XMPU_END_HI3 */
`define DDRMC5_NOC_XMPU_END_HI3_OFFSET 17'h12058
`define DDRMC5_NOC_XMPU_END_HI3_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI3_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI3_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI3_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI3_WIDTH 16

/* XMPU_MASTER3 */
`define DDRMC5_NOC_XMPU_MASTER3_OFFSET 17'h1205c
`define DDRMC5_NOC_XMPU_MASTER3_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER3_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER3_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER3_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER3_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER3_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER3_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER3_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER3_WIDTH 26

/* XMPU_CONFIG3 */
`define DDRMC5_NOC_XMPU_CONFIG3_OFFSET 17'h12060
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG3_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG3_WIDTH 5

/* XMPU_START_LO4 */
`define DDRMC5_NOC_XMPU_START_LO4_OFFSET 17'h12064
`define DDRMC5_NOC_XMPU_START_LO4_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO4_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO4_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO4_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO4_WIDTH 32

/* XMPU_START_HI4 */
`define DDRMC5_NOC_XMPU_START_HI4_OFFSET 17'h12068
`define DDRMC5_NOC_XMPU_START_HI4_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI4_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI4_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI4_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI4_WIDTH 16

/* XMPU_END_LO4 */
`define DDRMC5_NOC_XMPU_END_LO4_OFFSET 17'h1206c
`define DDRMC5_NOC_XMPU_END_LO4_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO4_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO4_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO4_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO4_WIDTH 32

/* XMPU_END_HI4 */
`define DDRMC5_NOC_XMPU_END_HI4_OFFSET 17'h12070
`define DDRMC5_NOC_XMPU_END_HI4_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI4_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI4_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI4_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI4_WIDTH 16

/* XMPU_MASTER4 */
`define DDRMC5_NOC_XMPU_MASTER4_OFFSET 17'h12074
`define DDRMC5_NOC_XMPU_MASTER4_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER4_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER4_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER4_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER4_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER4_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER4_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER4_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER4_WIDTH 26

/* XMPU_CONFIG4 */
`define DDRMC5_NOC_XMPU_CONFIG4_OFFSET 17'h12078
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG4_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG4_WIDTH 5

/* XMPU_START_LO5 */
`define DDRMC5_NOC_XMPU_START_LO5_OFFSET 17'h1207c
`define DDRMC5_NOC_XMPU_START_LO5_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO5_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO5_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO5_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO5_WIDTH 32

/* XMPU_START_HI5 */
`define DDRMC5_NOC_XMPU_START_HI5_OFFSET 17'h12080
`define DDRMC5_NOC_XMPU_START_HI5_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI5_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI5_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI5_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI5_WIDTH 16

/* XMPU_END_LO5 */
`define DDRMC5_NOC_XMPU_END_LO5_OFFSET 17'h12084
`define DDRMC5_NOC_XMPU_END_LO5_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO5_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO5_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO5_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO5_WIDTH 32

/* XMPU_END_HI5 */
`define DDRMC5_NOC_XMPU_END_HI5_OFFSET 17'h12088
`define DDRMC5_NOC_XMPU_END_HI5_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI5_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI5_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI5_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI5_WIDTH 16

/* XMPU_MASTER5 */
`define DDRMC5_NOC_XMPU_MASTER5_OFFSET 17'h1208c
`define DDRMC5_NOC_XMPU_MASTER5_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER5_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER5_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER5_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER5_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER5_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER5_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER5_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER5_WIDTH 26

/* XMPU_CONFIG5 */
`define DDRMC5_NOC_XMPU_CONFIG5_OFFSET 17'h12090
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG5_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG5_WIDTH 5

/* XMPU_START_LO6 */
`define DDRMC5_NOC_XMPU_START_LO6_OFFSET 17'h12094
`define DDRMC5_NOC_XMPU_START_LO6_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO6_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO6_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO6_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO6_WIDTH 32

/* XMPU_START_HI6 */
`define DDRMC5_NOC_XMPU_START_HI6_OFFSET 17'h12098
`define DDRMC5_NOC_XMPU_START_HI6_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI6_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI6_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI6_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI6_WIDTH 16

/* XMPU_END_LO6 */
`define DDRMC5_NOC_XMPU_END_LO6_OFFSET 17'h1209c
`define DDRMC5_NOC_XMPU_END_LO6_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO6_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO6_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO6_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO6_WIDTH 32

/* XMPU_END_HI6 */
`define DDRMC5_NOC_XMPU_END_HI6_OFFSET 17'h120a0
`define DDRMC5_NOC_XMPU_END_HI6_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI6_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI6_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI6_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI6_WIDTH 16

/* XMPU_MASTER6 */
`define DDRMC5_NOC_XMPU_MASTER6_OFFSET 17'h120a4
`define DDRMC5_NOC_XMPU_MASTER6_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER6_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER6_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER6_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER6_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER6_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER6_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER6_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER6_WIDTH 26

/* XMPU_CONFIG6 */
`define DDRMC5_NOC_XMPU_CONFIG6_OFFSET 17'h120a8
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG6_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG6_WIDTH 5

/* XMPU_START_LO7 */
`define DDRMC5_NOC_XMPU_START_LO7_OFFSET 17'h120ac
`define DDRMC5_NOC_XMPU_START_LO7_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO7_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO7_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO7_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO7_WIDTH 32

/* XMPU_START_HI7 */
`define DDRMC5_NOC_XMPU_START_HI7_OFFSET 17'h120b0
`define DDRMC5_NOC_XMPU_START_HI7_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI7_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI7_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI7_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI7_WIDTH 16

/* XMPU_END_LO7 */
`define DDRMC5_NOC_XMPU_END_LO7_OFFSET 17'h120b4
`define DDRMC5_NOC_XMPU_END_LO7_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO7_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO7_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO7_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO7_WIDTH 32

/* XMPU_END_HI7 */
`define DDRMC5_NOC_XMPU_END_HI7_OFFSET 17'h120b8
`define DDRMC5_NOC_XMPU_END_HI7_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI7_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI7_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI7_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI7_WIDTH 16

/* XMPU_MASTER7 */
`define DDRMC5_NOC_XMPU_MASTER7_OFFSET 17'h120bc
`define DDRMC5_NOC_XMPU_MASTER7_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER7_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER7_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER7_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER7_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER7_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER7_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER7_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER7_WIDTH 26

/* XMPU_CONFIG7 */
`define DDRMC5_NOC_XMPU_CONFIG7_OFFSET 17'h120c0
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG7_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG7_WIDTH 5

/* XMPU_START_LO8 */
`define DDRMC5_NOC_XMPU_START_LO8_OFFSET 17'h120c4
`define DDRMC5_NOC_XMPU_START_LO8_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO8_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO8_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO8_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO8_WIDTH 32

/* XMPU_START_HI8 */
`define DDRMC5_NOC_XMPU_START_HI8_OFFSET 17'h120c8
`define DDRMC5_NOC_XMPU_START_HI8_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI8_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI8_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI8_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI8_WIDTH 16

/* XMPU_END_LO8 */
`define DDRMC5_NOC_XMPU_END_LO8_OFFSET 17'h120cc
`define DDRMC5_NOC_XMPU_END_LO8_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO8_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO8_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO8_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO8_WIDTH 32

/* XMPU_END_HI8 */
`define DDRMC5_NOC_XMPU_END_HI8_OFFSET 17'h120d0
`define DDRMC5_NOC_XMPU_END_HI8_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI8_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI8_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI8_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI8_WIDTH 16

/* XMPU_MASTER8 */
`define DDRMC5_NOC_XMPU_MASTER8_OFFSET 17'h120d4
`define DDRMC5_NOC_XMPU_MASTER8_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER8_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER8_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER8_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER8_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER8_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER8_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER8_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER8_WIDTH 26

/* XMPU_CONFIG8 */
`define DDRMC5_NOC_XMPU_CONFIG8_OFFSET 17'h120d8
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG8_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG8_WIDTH 5

/* XMPU_START_LO9 */
`define DDRMC5_NOC_XMPU_START_LO9_OFFSET 17'h120dc
`define DDRMC5_NOC_XMPU_START_LO9_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO9_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO9_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO9_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO9_WIDTH 32

/* XMPU_START_HI9 */
`define DDRMC5_NOC_XMPU_START_HI9_OFFSET 17'h120e0
`define DDRMC5_NOC_XMPU_START_HI9_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI9_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI9_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI9_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI9_WIDTH 16

/* XMPU_END_LO9 */
`define DDRMC5_NOC_XMPU_END_LO9_OFFSET 17'h120e4
`define DDRMC5_NOC_XMPU_END_LO9_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO9_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO9_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO9_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO9_WIDTH 32

/* XMPU_END_HI9 */
`define DDRMC5_NOC_XMPU_END_HI9_OFFSET 17'h120e8
`define DDRMC5_NOC_XMPU_END_HI9_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI9_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI9_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI9_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI9_WIDTH 16

/* XMPU_MASTER9 */
`define DDRMC5_NOC_XMPU_MASTER9_OFFSET 17'h120ec
`define DDRMC5_NOC_XMPU_MASTER9_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER9_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER9_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER9_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER9_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER9_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER9_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER9_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER9_WIDTH 26

/* XMPU_CONFIG9 */
`define DDRMC5_NOC_XMPU_CONFIG9_OFFSET 17'h120f0
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG9_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG9_WIDTH 5

/* XMPU_START_LO10 */
`define DDRMC5_NOC_XMPU_START_LO10_OFFSET 17'h120f4
`define DDRMC5_NOC_XMPU_START_LO10_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO10_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO10_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO10_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO10_WIDTH 32

/* XMPU_START_HI10 */
`define DDRMC5_NOC_XMPU_START_HI10_OFFSET 17'h120f8
`define DDRMC5_NOC_XMPU_START_HI10_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI10_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI10_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI10_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI10_WIDTH 16

/* XMPU_END_LO10 */
`define DDRMC5_NOC_XMPU_END_LO10_OFFSET 17'h120fc
`define DDRMC5_NOC_XMPU_END_LO10_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO10_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO10_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO10_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO10_WIDTH 32

/* XMPU_END_HI10 */
`define DDRMC5_NOC_XMPU_END_HI10_OFFSET 17'h12100
`define DDRMC5_NOC_XMPU_END_HI10_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI10_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI10_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI10_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI10_WIDTH 16

/* XMPU_MASTER10 */
`define DDRMC5_NOC_XMPU_MASTER10_OFFSET 17'h12104
`define DDRMC5_NOC_XMPU_MASTER10_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER10_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER10_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER10_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER10_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER10_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER10_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER10_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER10_WIDTH 26

/* XMPU_CONFIG10 */
`define DDRMC5_NOC_XMPU_CONFIG10_OFFSET 17'h12108
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG10_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG10_WIDTH 5

/* XMPU_START_LO11 */
`define DDRMC5_NOC_XMPU_START_LO11_OFFSET 17'h1210c
`define DDRMC5_NOC_XMPU_START_LO11_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO11_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO11_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO11_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO11_WIDTH 32

/* XMPU_START_HI11 */
`define DDRMC5_NOC_XMPU_START_HI11_OFFSET 17'h12110
`define DDRMC5_NOC_XMPU_START_HI11_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI11_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI11_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI11_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI11_WIDTH 16

/* XMPU_END_LO11 */
`define DDRMC5_NOC_XMPU_END_LO11_OFFSET 17'h12114
`define DDRMC5_NOC_XMPU_END_LO11_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO11_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO11_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO11_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO11_WIDTH 32

/* XMPU_END_HI11 */
`define DDRMC5_NOC_XMPU_END_HI11_OFFSET 17'h12118
`define DDRMC5_NOC_XMPU_END_HI11_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI11_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI11_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI11_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI11_WIDTH 16

/* XMPU_MASTER11 */
`define DDRMC5_NOC_XMPU_MASTER11_OFFSET 17'h1211c
`define DDRMC5_NOC_XMPU_MASTER11_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER11_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER11_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER11_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER11_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER11_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER11_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER11_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER11_WIDTH 26

/* XMPU_CONFIG11 */
`define DDRMC5_NOC_XMPU_CONFIG11_OFFSET 17'h12120
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG11_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG11_WIDTH 5

/* XMPU_START_LO12 */
`define DDRMC5_NOC_XMPU_START_LO12_OFFSET 17'h12124
`define DDRMC5_NOC_XMPU_START_LO12_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO12_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO12_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO12_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO12_WIDTH 32

/* XMPU_START_HI12 */
`define DDRMC5_NOC_XMPU_START_HI12_OFFSET 17'h12128
`define DDRMC5_NOC_XMPU_START_HI12_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI12_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI12_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI12_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI12_WIDTH 16

/* XMPU_END_LO12 */
`define DDRMC5_NOC_XMPU_END_LO12_OFFSET 17'h1212c
`define DDRMC5_NOC_XMPU_END_LO12_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO12_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO12_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO12_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO12_WIDTH 32

/* XMPU_END_HI12 */
`define DDRMC5_NOC_XMPU_END_HI12_OFFSET 17'h12130
`define DDRMC5_NOC_XMPU_END_HI12_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI12_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI12_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI12_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI12_WIDTH 16

/* XMPU_MASTER12 */
`define DDRMC5_NOC_XMPU_MASTER12_OFFSET 17'h12134
`define DDRMC5_NOC_XMPU_MASTER12_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER12_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER12_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER12_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER12_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER12_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER12_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER12_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER12_WIDTH 26

/* XMPU_CONFIG12 */
`define DDRMC5_NOC_XMPU_CONFIG12_OFFSET 17'h12138
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG12_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG12_WIDTH 5

/* XMPU_START_LO13 */
`define DDRMC5_NOC_XMPU_START_LO13_OFFSET 17'h1213c
`define DDRMC5_NOC_XMPU_START_LO13_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO13_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO13_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO13_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO13_WIDTH 32

/* XMPU_START_HI13 */
`define DDRMC5_NOC_XMPU_START_HI13_OFFSET 17'h12140
`define DDRMC5_NOC_XMPU_START_HI13_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI13_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI13_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI13_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI13_WIDTH 16

/* XMPU_END_LO13 */
`define DDRMC5_NOC_XMPU_END_LO13_OFFSET 17'h12144
`define DDRMC5_NOC_XMPU_END_LO13_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO13_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO13_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO13_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO13_WIDTH 32

/* XMPU_END_HI13 */
`define DDRMC5_NOC_XMPU_END_HI13_OFFSET 17'h12148
`define DDRMC5_NOC_XMPU_END_HI13_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI13_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI13_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI13_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI13_WIDTH 16

/* XMPU_MASTER13 */
`define DDRMC5_NOC_XMPU_MASTER13_OFFSET 17'h1214c
`define DDRMC5_NOC_XMPU_MASTER13_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER13_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER13_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER13_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER13_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER13_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER13_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER13_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER13_WIDTH 26

/* XMPU_CONFIG13 */
`define DDRMC5_NOC_XMPU_CONFIG13_OFFSET 17'h12150
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG13_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG13_WIDTH 5

/* XMPU_START_LO14 */
`define DDRMC5_NOC_XMPU_START_LO14_OFFSET 17'h12154
`define DDRMC5_NOC_XMPU_START_LO14_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO14_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO14_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO14_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO14_WIDTH 32

/* XMPU_START_HI14 */
`define DDRMC5_NOC_XMPU_START_HI14_OFFSET 17'h12158
`define DDRMC5_NOC_XMPU_START_HI14_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI14_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI14_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI14_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI14_WIDTH 16

/* XMPU_END_LO14 */
`define DDRMC5_NOC_XMPU_END_LO14_OFFSET 17'h1215c
`define DDRMC5_NOC_XMPU_END_LO14_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO14_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO14_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO14_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO14_WIDTH 32

/* XMPU_END_HI14 */
`define DDRMC5_NOC_XMPU_END_HI14_OFFSET 17'h12160
`define DDRMC5_NOC_XMPU_END_HI14_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI14_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI14_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI14_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI14_WIDTH 16

/* XMPU_MASTER14 */
`define DDRMC5_NOC_XMPU_MASTER14_OFFSET 17'h12164
`define DDRMC5_NOC_XMPU_MASTER14_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER14_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER14_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER14_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER14_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER14_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER14_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER14_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER14_WIDTH 26

/* XMPU_CONFIG14 */
`define DDRMC5_NOC_XMPU_CONFIG14_OFFSET 17'h12168
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG14_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG14_WIDTH 5

/* XMPU_START_LO15 */
`define DDRMC5_NOC_XMPU_START_LO15_OFFSET 17'h1216c
`define DDRMC5_NOC_XMPU_START_LO15_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_START_LO15_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_START_LO15_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_START_LO15_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_START_LO15_WIDTH 32

/* XMPU_START_HI15 */
`define DDRMC5_NOC_XMPU_START_HI15_OFFSET 17'h12170
`define DDRMC5_NOC_XMPU_START_HI15_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_START_HI15_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI15_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_START_HI15_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_START_HI15_WIDTH 16

/* XMPU_END_LO15 */
`define DDRMC5_NOC_XMPU_END_LO15_OFFSET 17'h12174
`define DDRMC5_NOC_XMPU_END_LO15_FLD_RESERVED 11:0
`define DDRMC5_NOC_XMPU_END_LO15_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_XMPU_END_LO15_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_XMPU_END_LO15_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_XMPU_END_LO15_WIDTH 32

/* XMPU_END_HI15 */
`define DDRMC5_NOC_XMPU_END_HI15_OFFSET 17'h12178
`define DDRMC5_NOC_XMPU_END_HI15_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_XMPU_END_HI15_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI15_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_END_HI15_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_END_HI15_WIDTH 16

/* XMPU_MASTER15 */
`define DDRMC5_NOC_XMPU_MASTER15_OFFSET 17'h1217c
`define DDRMC5_NOC_XMPU_MASTER15_FLD_ID 9:0
`define DDRMC5_NOC_XMPU_MASTER15_FLD_ID_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER15_FLD_RESERVED 15:10
`define DDRMC5_NOC_XMPU_MASTER15_FLD_RESERVED_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER15_FLD_MASK 25:16
`define DDRMC5_NOC_XMPU_MASTER15_FLD_MASK_WIDTH 10
`define DDRMC5_NOC_XMPU_MASTER15_FLD_RESERVED_1 31:26
`define DDRMC5_NOC_XMPU_MASTER15_FLD_RESERVED_1_WIDTH 6
`define DDRMC5_NOC_XMPU_MASTER15_WIDTH 26

/* XMPU_CONFIG15 */
`define DDRMC5_NOC_XMPU_CONFIG15_OFFSET 17'h12180
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_ENABLE 0
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_ENABLE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_RDALLOWED 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_RDALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_WRALLOWED 2
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_WRALLOWED_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_REGIONNS 3
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_REGIONNS_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_NSCHECKTYPE 4
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_NSCHECKTYPE_WIDTH 1
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_RESERVED 31:5
`define DDRMC5_NOC_XMPU_CONFIG15_FLD_RESERVED_WIDTH 27
`define DDRMC5_NOC_XMPU_CONFIG15_WIDTH 5

/* REG_ADEC_CHK0 */
`define DDRMC5_NOC_REG_ADEC_CHK0_OFFSET 17'h12184
`define DDRMC5_NOC_REG_ADEC_CHK0_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_REG_ADEC_CHK0_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_REG_ADEC_CHK0_FLD_RESERVED 31:16
`define DDRMC5_NOC_REG_ADEC_CHK0_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_REG_ADEC_CHK0_WIDTH 16

/* REG_ADEC_CHK1 */
`define DDRMC5_NOC_REG_ADEC_CHK1_OFFSET 17'h12188
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_ENABLE 1:0
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_ENABLE_WIDTH 2
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_RESERVED 11:2
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_RESERVED_WIDTH 10
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_REG_ADEC_CHK1_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_REG_ADEC_CHK1_WIDTH 32

/* REG_ADEC_CHK2 */
`define DDRMC5_NOC_REG_ADEC_CHK2_OFFSET 17'h1218c
`define DDRMC5_NOC_REG_ADEC_CHK2_FLD_ADDR_HI 15:0
`define DDRMC5_NOC_REG_ADEC_CHK2_FLD_ADDR_HI_WIDTH 16
`define DDRMC5_NOC_REG_ADEC_CHK2_FLD_RESERVED 31:16
`define DDRMC5_NOC_REG_ADEC_CHK2_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_REG_ADEC_CHK2_WIDTH 16

/* REG_ADEC_CHK3 */
`define DDRMC5_NOC_REG_ADEC_CHK3_OFFSET 17'h12190
`define DDRMC5_NOC_REG_ADEC_CHK3_FLD_RESERVED 11:0
`define DDRMC5_NOC_REG_ADEC_CHK3_FLD_RESERVED_WIDTH 12
`define DDRMC5_NOC_REG_ADEC_CHK3_FLD_ADDR_LO 31:12
`define DDRMC5_NOC_REG_ADEC_CHK3_FLD_ADDR_LO_WIDTH 20
`define DDRMC5_NOC_REG_ADEC_CHK3_WIDTH 32

/* XMPU_LOCK */
`define DDRMC5_NOC_XMPU_LOCK_OFFSET 17'h12194
`define DDRMC5_NOC_XMPU_LOCK_FLD_PROT 0
`define DDRMC5_NOC_XMPU_LOCK_FLD_PROT_WIDTH 1
`define DDRMC5_NOC_XMPU_LOCK_WIDTH 1

/* ADEC_LOCK */
`define DDRMC5_NOC_ADEC_LOCK_OFFSET 17'h12198
`define DDRMC5_NOC_ADEC_LOCK_FLD_PROT 0
`define DDRMC5_NOC_ADEC_LOCK_FLD_PROT_WIDTH 1
`define DDRMC5_NOC_ADEC_LOCK_WIDTH 1

/* XMPU_ERR_STATUS */
`define DDRMC5_NOC_XMPU_ERR_STATUS_OFFSET 17'h1219c
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RESERVED 0
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RDPERMVIO 1
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RDPERMVIO_WIDTH 1
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_WRPERMVIO 2
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_WRPERMVIO_WIDTH 1
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_SECURITYVIO 3
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_SECURITYVIO_WIDTH 1
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_REGIONVIO 8:4
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_REGIONVIO_WIDTH 5
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RESERVED_1 31:9
`define DDRMC5_NOC_XMPU_ERR_STATUS_FLD_RESERVED_1_WIDTH 23
`define DDRMC5_NOC_XMPU_ERR_STATUS_WIDTH 9

/* XMPU_ERR_ADD_LO0 */
`define DDRMC5_NOC_XMPU_ERR_ADD_LO0_OFFSET 17'h121a0
`define DDRMC5_NOC_XMPU_ERR_ADD_LO0_FLD_XMPU_ERR_ADD_LO 31:0
`define DDRMC5_NOC_XMPU_ERR_ADD_LO0_FLD_XMPU_ERR_ADD_LO_WIDTH 32
`define DDRMC5_NOC_XMPU_ERR_ADD_LO0_WIDTH 32

/* XMPU_ERR_ADD_HI0 */
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_OFFSET 17'h121a4
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_FLD_XMPU_ERR_ADD_HI 15:0
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_FLD_XMPU_ERR_ADD_HI_WIDTH 16
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_FLD_RESERVED 31:16
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_FLD_RESERVED_WIDTH 16
`define DDRMC5_NOC_XMPU_ERR_ADD_HI0_WIDTH 16

/* XMPU_ERR_AXI_ID */
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_OFFSET 17'h121a8
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_FLD_XMPU_ERR_SMID 9:0
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_FLD_XMPU_ERR_SMID_WIDTH 10
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_FLD_RESERVED 31:10
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_FLD_RESERVED_WIDTH 22
`define DDRMC5_NOC_XMPU_ERR_AXI_ID_WIDTH 10

/* ADEC_CHK_ERR_LOG */
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_OFFSET 17'h121ac
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_LT_LOW_REGION_VIO 0
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_LT_LOW_REGION_VIO_WIDTH 1
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_GT_LOW_REGION_VIO 1
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_GT_LOW_REGION_VIO_WIDTH 1
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_LT_HIGH_REGION_VIO 2
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_LT_HIGH_REGION_VIO_WIDTH 1
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_GT_HIGH_REGION_VIO 3
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_GT_HIGH_REGION_VIO_WIDTH 1
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_RESERVED 31:4
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_FLD_RESERVED_WIDTH 28
`define DDRMC5_NOC_ADEC_CHK_ERR_LOG_WIDTH 4

/* REG_ADEC17 */
`define DDRMC5_NOC_REG_ADEC17_OFFSET 17'h121b0
`define DDRMC5_NOC_REG_ADEC17_FLD_ROW_MASK 17:0
`define DDRMC5_NOC_REG_ADEC17_FLD_ROW_MASK_WIDTH 18
`define DDRMC5_NOC_REG_ADEC17_FLD_COL_MASK 28:18
`define DDRMC5_NOC_REG_ADEC17_FLD_COL_MASK_WIDTH 11
`define DDRMC5_NOC_REG_ADEC17_FLD_BANK_MASK 30:29
`define DDRMC5_NOC_REG_ADEC17_FLD_BANK_MASK_WIDTH 2
`define DDRMC5_NOC_REG_ADEC17_FLD_RESERVED 31
`define DDRMC5_NOC_REG_ADEC17_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_ADEC17_WIDTH 31

/* REG_ADEC18 */
`define DDRMC5_NOC_REG_ADEC18_OFFSET 17'h121b4
`define DDRMC5_NOC_REG_ADEC18_FLD_RANK_MASK 1:0
`define DDRMC5_NOC_REG_ADEC18_FLD_RANK_MASK_WIDTH 2
`define DDRMC5_NOC_REG_ADEC18_FLD_LRANK_MASK 5:2
`define DDRMC5_NOC_REG_ADEC18_FLD_LRANK_MASK_WIDTH 4
`define DDRMC5_NOC_REG_ADEC18_FLD_CH_MASK 6
`define DDRMC5_NOC_REG_ADEC18_FLD_CH_MASK_WIDTH 1
`define DDRMC5_NOC_REG_ADEC18_FLD_GROUP_MASK 9:7
`define DDRMC5_NOC_REG_ADEC18_FLD_GROUP_MASK_WIDTH 3
`define DDRMC5_NOC_REG_ADEC18_FLD_RESERVED 31:10
`define DDRMC5_NOC_REG_ADEC18_FLD_RESERVED_WIDTH 22
`define DDRMC5_NOC_REG_ADEC18_WIDTH 10

/* REG_ADEC19 */
`define DDRMC5_NOC_REG_ADEC19_OFFSET 17'h121b8
`define DDRMC5_NOC_REG_ADEC19_FLD_ROW_MATCH 17:0
`define DDRMC5_NOC_REG_ADEC19_FLD_ROW_MATCH_WIDTH 18
`define DDRMC5_NOC_REG_ADEC19_FLD_COL_MATCH 28:18
`define DDRMC5_NOC_REG_ADEC19_FLD_COL_MATCH_WIDTH 11
`define DDRMC5_NOC_REG_ADEC19_FLD_BANK_MATCH 30:29
`define DDRMC5_NOC_REG_ADEC19_FLD_BANK_MATCH_WIDTH 2
`define DDRMC5_NOC_REG_ADEC19_FLD_RESERVED 31
`define DDRMC5_NOC_REG_ADEC19_FLD_RESERVED_WIDTH 1
`define DDRMC5_NOC_REG_ADEC19_WIDTH 31

/* REG_ADEC20 */
`define DDRMC5_NOC_REG_ADEC20_OFFSET 17'h121bc
`define DDRMC5_NOC_REG_ADEC20_FLD_RANK_MATCH 1:0
`define DDRMC5_NOC_REG_ADEC20_FLD_RANK_MATCH_WIDTH 2
`define DDRMC5_NOC_REG_ADEC20_FLD_LRANK_MATCH 5:2
`define DDRMC5_NOC_REG_ADEC20_FLD_LRANK_MATCH_WIDTH 4
`define DDRMC5_NOC_REG_ADEC20_FLD_CH_MATCH 6
`define DDRMC5_NOC_REG_ADEC20_FLD_CH_MATCH_WIDTH 1
`define DDRMC5_NOC_REG_ADEC20_FLD_PERSISTENT 7
`define DDRMC5_NOC_REG_ADEC20_FLD_PERSISTENT_WIDTH 1
`define DDRMC5_NOC_REG_ADEC20_FLD_DONE 8
`define DDRMC5_NOC_REG_ADEC20_FLD_DONE_WIDTH 1
`define DDRMC5_NOC_REG_ADEC20_FLD_MATCH_EN 9
`define DDRMC5_NOC_REG_ADEC20_FLD_MATCH_EN_WIDTH 1
`define DDRMC5_NOC_REG_ADEC20_FLD_GROUP_MATCH 12:10
`define DDRMC5_NOC_REG_ADEC20_FLD_GROUP_MATCH_WIDTH 3
`define DDRMC5_NOC_REG_ADEC20_FLD_RESERVED 31:13
`define DDRMC5_NOC_REG_ADEC20_FLD_RESERVED_WIDTH 19
`define DDRMC5_NOC_REG_ADEC20_WIDTH 13

/* REG_ADEC21 */
`define DDRMC5_NOC_REG_ADEC21_OFFSET 17'h121c0
`define DDRMC5_NOC_REG_ADEC21_FLD_DONE_CRYPTO 0
`define DDRMC5_NOC_REG_ADEC21_FLD_DONE_CRYPTO_WIDTH 1
`define DDRMC5_NOC_REG_ADEC21_FLD_MATCH_EN_CRYPTO 1
`define DDRMC5_NOC_REG_ADEC21_FLD_MATCH_EN_CRYPTO_WIDTH 1
`define DDRMC5_NOC_REG_ADEC21_FLD_RESERVED 31:2
`define DDRMC5_NOC_REG_ADEC21_FLD_RESERVED_WIDTH 30
`define DDRMC5_NOC_REG_ADEC21_WIDTH 2

/* ADD_PAR_ERR_INJ_ADEC */
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_OFFSET 17'h121c4
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_EN0 0
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_EN0_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_PERSISTENT0 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_PERSISTENT0_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADDRESS_TYPE0 3:2
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADDRESS_TYPE0_WIDTH 2
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_DONE0 4
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_DONE0_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_DRAM_RANK0 6:5
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_DRAM_RANK0_WIDTH 2
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_EN1 7
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_EN1_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_PERSISTENT1 8
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_PERSISTENT1_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADDRESS_TYPE1 10:9
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADDRESS_TYPE1_WIDTH 2
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_DONE1 11
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ERR_INJ_DONE1_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_DRAM_RANK1 13:12
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_DRAM_RANK1_WIDTH 2
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_CHK_EN0 14
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_CHK_EN0_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_LOG_EN0 15
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_LOG_EN0_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_CHK_EN1 16
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_CHK_EN1_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_LOG_EN1 17
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_ADEC_ADDR_PAR_LOG_EN1_WIDTH 1
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_RESERVED 31:18
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_FLD_RESERVED_WIDTH 14
`define DDRMC5_NOC_ADD_PAR_ERR_INJ_ADEC_WIDTH 18

/* ADEC_ADD_PAR_ERR_LOG0_0 */
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_0_OFFSET 17'h121c8
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_0_WIDTH 32

/* ADEC_ADD_PAR_ERR_LOG1_0 */
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_0_OFFSET 17'h121cc
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_0_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_0_WIDTH 32

/* ADEC_ADD_PAR_ERR_LOG0_1 */
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_1_OFFSET 17'h121d0
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG0_1_WIDTH 32

/* ADEC_ADD_PAR_ERR_LOG1_1 */
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_1_OFFSET 17'h121d4
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO 31:0
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_1_FLD_ERR_LOG_INFO_WIDTH 32
`define DDRMC5_NOC_ADEC_ADD_PAR_ERR_LOG1_1_WIDTH 32

// spyglass enable_block ConstName

`endif
