
//------> /softs/mentor/cpult/10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /softs/mentor/cpult/10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   dirren@lapsrv6.epfl.ch
//  Generated date: Wed Mar  8 15:22:31 2023
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    main_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module main_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for main_core_core_fsm_1
  parameter
    core_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : main_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    main_core
// ------------------------------------------------------------------


module main_core (
  clk, rst, return_rsc_dat, return_rsc_triosy_lz
);
  input clk;
  input rst;
  output [31:0] return_rsc_dat;
  output return_rsc_triosy_lz;


  // Interconnect Declarations
  reg return_rsc_triosy_obj_ld;
  wire [2:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_v1 #(.rscid(32'sd4),
  .width(32'sd32)) return_rsci (
      .idat(32'b00000000000000000000000000000001),
      .dat(return_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_rsc_triosy_obj (
      .ld(return_rsc_triosy_obj_ld),
      .lz(return_rsc_triosy_lz)
    );
  main_core_core_fsm main_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  always @(posedge clk) begin
    if ( rst ) begin
      return_rsc_triosy_obj_ld <= 1'b0;
    end
    else begin
      return_rsc_triosy_obj_ld <= ~ (fsm_output[1]);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    main
// ------------------------------------------------------------------


module main (
  clk, rst, return_rsc_dat, return_rsc_triosy_lz
);
  input clk;
  input rst;
  output [31:0] return_rsc_dat;
  output return_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  main_core main_core_inst (
      .clk(clk),
      .rst(rst),
      .return_rsc_dat(return_rsc_dat),
      .return_rsc_triosy_lz(return_rsc_triosy_lz)
    );
endmodule



