// tb.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module tb (
	);

	wire         clock_reset_inst_clock_clk;                                                     // clock_reset_inst:clock -> [component_dpi_controller_example_inst:clock, example_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                   // clock_reset_inst:clock2x -> [component_dpi_controller_example_inst:clock2x, main_dpi_controller_inst:clock2x]
	wire         component_dpi_controller_example_inst_component_call_valid;                     // component_dpi_controller_example_inst:start -> example_inst:start
	wire         example_inst_call_stall;                                                        // example_inst:busy -> component_dpi_controller_example_inst:busy
	wire         component_dpi_controller_example_inst_component_done_conduit;                   // component_dpi_controller_example_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                             // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_example_inst_component_wait_for_stream_writes_conduit; // component_dpi_controller_example_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         component_dpi_controller_example_inst_dpi_control_bind_conduit;                 // component_dpi_controller_example_inst:bind_interfaces -> example_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_example_inst_dpi_control_enable_conduit;               // component_dpi_controller_example_inst:enable_interfaces -> example_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         concatenate_component_done_inst_out_conduit_conduit;                            // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;          // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         split_component_start_inst_out_conduit_0_conduit;                               // split_component_start_inst:out_conduit_0 -> component_dpi_controller_example_inst:component_enabled
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                    // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         example_inst_return_valid;                                                      // example_inst:done -> component_dpi_controller_example_inst:done
	wire         component_dpi_controller_example_inst_component_return_stall;                   // component_dpi_controller_example_inst:stall -> example_inst:stall
	wire  [31:0] example_inst_returndata_data;                                                   // example_inst:returndata -> component_dpi_controller_example_inst:returndata
	wire         clock_reset_inst_reset_reset;                                                   // clock_reset_inst:resetn -> [component_dpi_controller_example_inst:resetn, example_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn]
	wire         component_dpi_controller_example_inst_component_irq_irq;                        // irq_mapper:sender_irq -> component_dpi_controller_example_inst:done_irq

	clock_reset clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //  output,  width = 1,      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //  output,  width = 1,      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //  output,  width = 1,    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  //   input,  width = 1, reset_ctrl.conduit
	);

	dpic_example component_dpi_controller_example_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                     //   input,   width = 1,                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                   //   input,   width = 1,                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                   //   input,   width = 1,                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_example_inst_dpi_control_bind_conduit),                 //  output,   width = 1,                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_example_inst_dpi_control_enable_conduit),               //  output,   width = 1,               dpi_control_enable.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                               //   input,   width = 1,                component_enabled.conduit
		.component_done                   (component_dpi_controller_example_inst_component_done_conduit),                   //  output,   width = 1,                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_example_inst_component_wait_for_stream_writes_conduit), //  output,   width = 1, component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                               //   input,   width = 1,                       agent_busy.conduit
		.read_implicit_streams            (),                                                                               //  output,   width = 1,            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                               //  output,   width = 1,             readback_from_agents.conduit
		.start                            (component_dpi_controller_example_inst_component_call_valid),                     //  output,   width = 1,                   component_call.valid
		.busy                             (example_inst_call_stall),                                                        //   input,   width = 1,                                 .stall
		.done                             (example_inst_return_valid),                                                      //   input,   width = 1,                 component_return.valid
		.stall                            (component_dpi_controller_example_inst_component_return_stall),                   //  output,   width = 1,                                 .stall
		.done_irq                         (component_dpi_controller_example_inst_component_irq_irq),                        //   input,   width = 1,                    component_irq.irq
		.returndata                       (example_inst_returndata_data)                                                    //   input,  width = 32,                       returndata.data
	);

	cat_done concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),          //  output,  width = 1,  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_example_inst_component_done_conduit)  //   input,  width = 1, in_conduit_0.conduit
	);

	cat_cwfsw concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),          //  output,  width = 1,  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_example_inst_component_wait_for_stream_writes_conduit)  //   input,  width = 1, in_conduit_0.conduit
	);

	example_cfan example_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit (component_dpi_controller_example_inst_dpi_control_bind_conduit)  //   input,  width = 1, in_conduit.conduit
	);

	example_en_cfan example_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit (component_dpi_controller_example_inst_dpi_control_enable_conduit)  //   input,  width = 1, in_conduit.conduit
	);

	example example_inst (
		.clock      (clock_reset_inst_clock_clk),                                   //   input,   width = 1,      clock.clk
		.resetn     (clock_reset_inst_reset_reset),                                 //   input,   width = 1,      reset.reset_n
		.start      (component_dpi_controller_example_inst_component_call_valid),   //   input,   width = 1,       call.valid
		.busy       (example_inst_call_stall),                                      //  output,   width = 1,           .stall
		.done       (example_inst_return_valid),                                    //  output,   width = 1,     return.valid
		.stall      (component_dpi_controller_example_inst_component_return_stall), //   input,   width = 1,           .stall
		.returndata (example_inst_returndata_data)                                  //  output,  width = 32, returndata.data
	);

	main_dpi_controller main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //   input,  width = 1,                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //   input,  width = 1,                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //   input,  width = 1,                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //  output,  width = 1,                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //   input,  width = 1,                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), //   input,  width = 1, component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //  output,  width = 1,                       reset_ctrl.conduit
	);

	sp_cstart split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //   input,  width = 1,    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    //  output,  width = 1, out_conduit_0.conduit
	);

	tb_altera_irq_mapper_1920_trjgw7i irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                              //   input,  width = 1,       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                           //   input,  width = 1, clk_reset.reset
		.sender_irq (component_dpi_controller_example_inst_component_irq_irq)  //  output,  width = 1,    sender.irq
	);

endmodule
