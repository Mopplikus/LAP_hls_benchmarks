// tb_kernel_3mm_inst.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module tb_kernel_3mm_inst (
		input  wire [63:0] A,                    //         A.data
		input  wire [63:0] B,                    //         B.data
		input  wire [63:0] C,                    //         C.data
		input  wire [63:0] D,                    //         D.data
		input  wire [63:0] E,                    //         E.data
		input  wire [63:0] F,                    //         F.data
		input  wire [63:0] G,                    //         G.data
		output wire [31:0] avmm_1_rw_address,    // avmm_1_rw.address
		output wire [3:0]  avmm_1_rw_byteenable, //          .byteenable
		output wire        avmm_1_rw_read,       //          .read
		input  wire [31:0] avmm_1_rw_readdata,   //          .readdata
		output wire        avmm_1_rw_write,      //          .write
		output wire [31:0] avmm_1_rw_writedata,  //          .writedata
		input  wire        start,                //      call.valid
		output wire        busy,                 //          .stall
		input  wire        clock,                //     clock.clk
		input  wire        resetn,               //     reset.reset_n
		output wire        done,                 //    return.valid
		input  wire        stall                 //          .stall
	);

	kernel_3mm_internal kernel_3mm_internal_inst (
		.clock                (clock),                //     clock.clk
		.resetn               (resetn),               //     reset.reset_n
		.start                (start),                //      call.valid
		.busy                 (busy),                 //          .stall
		.done                 (done),                 //    return.valid
		.stall                (stall),                //          .stall
		.A                    (A),                    //         A.data
		.B                    (B),                    //         B.data
		.C                    (C),                    //         C.data
		.D                    (D),                    //         D.data
		.E                    (E),                    //         E.data
		.F                    (F),                    //         F.data
		.G                    (G),                    //         G.data
		.avmm_1_rw_address    (avmm_1_rw_address),    // avmm_1_rw.address
		.avmm_1_rw_byteenable (avmm_1_rw_byteenable), //          .byteenable
		.avmm_1_rw_read       (avmm_1_rw_read),       //          .read
		.avmm_1_rw_readdata   (avmm_1_rw_readdata),   //          .readdata
		.avmm_1_rw_write      (avmm_1_rw_write),      //          .write
		.avmm_1_rw_writedata  (avmm_1_rw_writedata)   //          .writedata
	);

endmodule
