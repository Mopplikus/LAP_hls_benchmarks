// matvec.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module matvec (
		input  wire        clock,  //  clock.clk
		input  wire        resetn, //  reset.reset_n
		input  wire        start,  //   call.valid
		output wire        busy,   //       .stall
		output wire        done,   // return.valid
		input  wire        stall,  //       .stall
		input  wire [63:0] M,      //      M.data
		input  wire [63:0] V,      //      V.data
		input  wire [63:0] Out0    //   Out0.data
	);

	matvec_internal matvec_internal_inst (
		.clock  (clock),  //   input,   width = 1,  clock.clk
		.resetn (resetn), //   input,   width = 1,  reset.reset_n
		.start  (start),  //   input,   width = 1,   call.valid
		.busy   (busy),   //  output,   width = 1,       .stall
		.done   (done),   //  output,   width = 1, return.valid
		.stall  (stall),  //   input,   width = 1,       .stall
		.M      (M),      //   input,  width = 64,      M.data
		.V      (V),      //   input,  width = 64,      V.data
		.Out0   (Out0)    //   input,  width = 64,   Out0.data
	);

endmodule
