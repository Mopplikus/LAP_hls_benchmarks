`ifndef _noc_ddrmc5_define_vh_
`define _noc_ddrmc5_define_vh_

`define D5_NOC_DDRMC5_RETURN_ID_WIDTH  2
`define D5_NOC_NPS_DDRMC5_VC           5

`endif
