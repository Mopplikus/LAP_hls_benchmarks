// triangular.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module triangular (
		input  wire        clock,  //  clock.clk
		input  wire        resetn, //  reset.reset_n
		input  wire        start,  //   call.valid
		output wire        busy,   //       .stall
		output wire        done,   // return.valid
		input  wire        stall,  //       .stall
		input  wire [63:0] x,      //      x.data
		input  wire [63:0] A,      //      A.data
		input  wire [31:0] n       //      n.data
	);

	triangular_internal triangular_internal_inst (
		.clock  (clock),  //   input,   width = 1,  clock.clk
		.resetn (resetn), //   input,   width = 1,  reset.reset_n
		.start  (start),  //   input,   width = 1,   call.valid
		.busy   (busy),   //  output,   width = 1,       .stall
		.done   (done),   //  output,   width = 1, return.valid
		.stall  (stall),  //   input,   width = 1,       .stall
		.x      (x),      //   input,  width = 64,      x.data
		.A      (A),      //   input,  width = 64,      A.data
		.n      (n)       //   input,  width = 32,      n.data
	);

endmodule
