    .INIT_00(256'h0148062b40f2002002f30c2b20f2ff00014308208ac01f000148083660728000),
    .INIT_01(256'h0149082f01f2075402f80d2262c0100101480801002200490149082b80f20033),
    .INIT_02(256'h0143081d0021d002001303220083205d0142062076a1d0010142000108220745),
    .INIT_03(256'h00b0021d0101d010001301326263226c02f20e1d0081d000014208326263214c),
    .INIT_04(256'h037000207421d00802f30f36618324f80043001d0201d0040140063262632433),
    .INIT_05(256'h02f20d2262c0106002f20c01002322330012ff207481d0820250000504032597),
    .INIT_06(256'h025000030bf20711037000207422075402f20f3661f0109f02f20e1d04020748),
    .INIT_07(256'h020c391d08022ffd00b1172262c206e300b01601002207290013002074820719),
    .INIT_08(256'h001301207480b00002f220030bf3202f02f117207420d08002f0163601709002),
    .INIT_09(256'h02f018208ac011ff020c3920134010ff00b1192262c3602f00b018010020d001),
    .INIT_0A(256'h00b01a010001b200001302207481b10002f221050401900102f119207420121f),
    .INIT_0B(256'h02f11b0900d0900102f01a220082f000020c39207820100100b11b207543e029),
    .INIT_0C(256'h00b11d0900d2b00000b01c25000250000013033662f3202f02f2220d0800d040),
    .INIT_0D(256'h02f223014d00900102f11d250002be0f02f01c366332bf7e020c390d0402b00c),
    .INIT_0E(256'h01f1ff1dedb0d02001d0ff0bf050900d0012000be042d001025000015090300f),
    .INIT_0F(256'h0140060144009006014006226412203a0140063263f090060310001ff323603f),
    .INIT_10(256'h0141000b014360460140060b2150d080014100013000900d0140060150a09006),
    .INIT_11(256'h0100300d0080900701400e143000900701400e142002204101400e0d01009007),
    .INIT_12(256'h022ffd011012071b022ffd030072070b025000143002072700b2241420025000),
    .INIT_13(256'h022ffd2264c20729022ffd1410620719022ffd3a6502072b022ffd19001206e7),
    .INIT_14(256'h022ffd2d2092072d022ffd2d30a206e7022ffd1235020703022ffd1024020725),
    .INIT_15(256'h022ffd01a00206e3022ffd25000206eb022ffd02010206e7022ffd09008206ed),
    .INIT_16(256'h022ffd09c1c3e05a022ffd14b0619001022ffd14b0601019022ffd0bb1325000),
    .INIT_17(256'h022ffd10ba0200e3022ffd09f1f200fd022ffd09e1e200f5022ffd09d1d25000),
    .INIT_18(256'h022ffd13f002089d022ffd13e0032060022ffd13d000d001022ffd10cb00900d),
    .INIT_19(256'h022ffd2062f208be022ffd20681208db022ffd01b0001101022ffd01a0401080),
    .INIT_1A(256'h022ffd2062f01000022ffd09d0736063022ffd2062f1dc93022ffd09c07208eb),
    .INIT_1B(256'h022ffd01aeb2f002022ffd09f0701000022ffd2062f2f001022ffd09e0705001),
    .INIT_1C(256'h022ffd0b6121d102022ffd0b5110311e022ffd0b410001e0022ffd01b0120b4d),
    .INIT_1D(256'h022ffd12e601d104022ffd12d5032082022ffd10c401d110022ffd0360132080),
    .INIT_1E(256'h022ffd3e6751d116022ffd1bb003208e022ffd19a011d112022ffd13f003208c),
    .INIT_1F(256'h022ffd2068122017022ffd01b0132087022ffd01aec1d100022ffd2500032094),
    .INIT_20(256'h022ffd2063301220022ffd2df07001d0022ffd20633320a8022ffd2500001200),
    .INIT_21(256'h022ffd20633001d0022ffd2dd0722094022ffd20633320a8022ffd2de071d190),
    .INIT_22(256'h022ffd2063322094022ffd2db07320a8022ffd206331d1b0022ffd2dc0701220),
    .INIT_23(256'h022ffd0150001204022ffd0146c001d0022ffd25000320a8022ffd2da0701203),
    .INIT_24(256'h022ffd0d010320a8022ffd0b0141d1b0022ffd0b215320a8022ffd013001d190),
    .INIT_25(256'h022ffd142000dd40022ffd0d0083609b022ffd143000dd10022ffd1420001000),
    .INIT_26(256'h022ffd190012f002022ffd0110114000022ffd030070dd20022ffd1430014000),
    .INIT_27(256'h022ffd10240320a4022ffd2269b1d112022ffd14106320a2022ffd3a69f1d110),
    .INIT_28(256'h022ffd09008320a8022ffd2d20901222022ffd2d30a320a6022ffd123501d116),
    .INIT_29(256'h022ffd2d008320a8022ffd2d20901226022ffd2d30a320a8022ffd0601001223),
    .INIT_2A(256'h022ffd14c002f03a022ffd14b0001000022ffd14a06200df022ffd250002f239),
    .INIT_2B(256'h022ffd250002f024022ffd14f0001001022ffd14e000d004022ffd14d0009002),
    .INIT_2C(256'h022ffd39000208a6022ffd190e9208a9022ffd3900020108022ffd110b9200ef),
    .INIT_2D(256'h022ffd390002b02e022ffd1100720914022ffd3e6ba2b02e022ffd19011208ac),
    .INIT_2E(256'h022ffd25000200e9022ffd1100a200df022ffd250002089d022ffd190f620914),
    .INIT_2F(256'h022ffd2073709001022ffd206ce2b04e022ffd206c4200df022ffd00c0020126),
    .INIT_30(256'h022ffd2500009002022ffd20737320d4022ffd206ce1d001022ffd206c40300f),
    .INIT_31(256'h022ffd14c062b20f022ffd14100208ac022ffd14c06320ce022ffd011000d002),
    .INIT_32(256'h022ffd14c0620754022ffd1410001002022ffd14c062b80f022ffd141002b40f),
    .INIT_33(256'h022ffd3a6d1208ac022ffd1d10a20134022ffd2500022008022ffd1410020782),
    .INIT_34(256'h022ffd01a0022008022ffd2500020782022ffd1113020754022ffd1110701000),
    .INIT_35(256'h022ffd390002b80f022ffd206b02b40f022ffd090062b20f022ffd2073a208ac),
    .INIT_36(256'h022ffd366d920709022ffd1910120770022ffd206a92f032022ffd0110401001),
    .INIT_37(256'h022ffd207372071f022ffd206ce22481022ffd00100206e5022ffd04a00206e9),
    .INIT_38(256'h022ffd0110d20713022ffd2500025000022ffd366d4206e3022ffd1920120717),
    .INIT_39(256'h022ffd0115f206e5022ffd2273720721022ffd0112020703022ffd2273720707),
    .INIT_3A(256'h022ffd0113120713022ffd227372071d022ffd0113e20713022ffd2273725000),
    .INIT_3B(256'h022ffd0113020725022ffd2273725000022ffd01133206e5022ffd2273720729),
    .INIT_3C(256'h022ffd01132206e5022ffd2273720717022ffd0113120705022ffd2273720709),
    .INIT_3D(256'h022ffd01134206e5022ffd2273720727022ffd011332070d022ffd2273725000),
    .INIT_3E(256'h022ffd01136206e3022ffd22737206bc022ffd011350300f022ffd2273709001),
    .INIT_3F(256'h022ffd01138206e5022ffd227372070d022ffd0113720703022ffd2273725000),
    .INIT_40(256'h022ffd011411400e022ffd227371400e022ffd0113903008022ffd2273709002),
    .INIT_41(256'h022ffd0114325000022ffd22737206e3022ffd01142206bc022ffd227371400e),
    .INIT_42(256'h022ffd0114501f00022ffd22737208db022ffd0114401100022ffd22737010c0),
    .INIT_43(256'h022ffd01147208f5022ffd2273701c00022ffd0114601d01022ffd2273701e00),
    .INIT_44(256'h022ffd0114901f00022ffd22737208db022ffd0114801100022ffd22737010a0),
    .INIT_45(256'h022ffd0114b208f5022ffd2273701c00022ffd0114a01d00022ffd2273701e00),
    .INIT_46(256'h022ffd0114d208f2022ffd22737208db022ffd0114c01101022ffd22737010c0),
    .INIT_47(256'h022ffd0114f03c3f022ffd2273703d7c022ffd0114e03e3c022ffd2273703f81),
    .INIT_48(256'h022ffd0115105c00022ffd2273705d03022ffd0115005e40022ffd2273705f00),
    .INIT_49(256'h022ffd0115301101022ffd22737010c0022ffd0115225000022ffd22737208f5),
    .INIT_4A(256'h022ffd0115503e7f022ffd2273703fff022ffd01154208f2022ffd22737208db),
    .INIT_4B(256'h022ffd0115705e80022ffd2273705f00022ffd0115603cff022ffd2273703dfd),
    .INIT_4C(256'h022ffd0115925000022ffd22737208f5022ffd0115805c00022ffd2273705d00),
    .INIT_4D(256'h022ffd2073e208f2022ffd22737208db022ffd0115a01101022ffd22737010c0),
    .INIT_4E(256'h022ffd0d02003cff022ffd0900d03dfe022ffd2500003eff022ffd2d10603fff),
    .INIT_4F(256'h022ffd0d01001101022ffd0900d010c0022ffd2500025000022ffd3673a208f5),
    .INIT_50(256'h022ffd0306003eff022ffd0900003fff022ffd25000208f2022ffd3673e208db),
    .INIT_51(256'h022ffd2500005e00022ffd0309f05f00022ffd0900003cff022ffd2500003dfe),
    .INIT_52(256'h022ffd0410025000022ffd20745208f5022ffd0316005c00022ffd0010005d01),
    .INIT_53(256'h022ffd206e50900f022ffd207072f01e022ffd2070d2f032022ffd2d10001000),
    .INIT_54(256'h022ffd2500036192022ffd206e30d020022ffd206bc36192022ffd207420d040),
    .INIT_55(256'h022ffd041000d080022ffd207420900e022ffd0319f3618d022ffd001000d080),
    .INIT_56(256'h022ffd206e50d020022ffd2070736186022ffd207270d040022ffd2d10036189),
    .INIT_57(256'h022ffd207450900e022ffd3277e36180022ffd1d0010d010022ffd0b03236183),
    .INIT_58(256'h022ffd207272f00b022ffd250000901b022ffd206e332169022ffd206bc0d004),
    .INIT_59(256'h022ffd206bc36176022ffd010021d0e0022ffd206e5030f0022ffd207072b04e),
    .INIT_5A(256'h022ffd0319f36176022ffd001000d020022ffd250000900d022ffd206e322177),
    .INIT_5B(256'h022ffd2500022177022ffd2d10036170022ffd041001d049022ffd2074209006),
    .INIT_5C(256'h022ffd2d103206e3022ffd0b13220727022ffd2076a36176022ffd010001d053),
    .INIT_5D(256'h022ffd0b03220713022ffd206e522008022ffd2070720782022ffd207272078b),
    .INIT_5E(256'h022ffd206bc208ac022ffd0104020134022ffd3277e2089d022ffd1d001206e3),
    .INIT_5F(256'h022ffd206bc22008022ffd0102020782022ffd2500020754022ffd206e301000),
    .INIT_60(256'h022ffd1d0002b20e022ffd2074522190022ffd2500001080022ffd206e32b10e),
    .INIT_61(256'h022ffd206e501020022ffd206e92b40e022ffd2071f22190022ffd3278901040),
    .INIT_62(256'h022ffd2072701010022ffd227862b80e022ffd207132089d022ffd2500022190),
    .INIT_63(256'h022ffd206bd01008022ffd0bc022b80f022ffd206e52089d022ffd2071d22190),
    .INIT_64(256'h022ffd207252b40f022ffd2074d2089d022ffd2075922209022ffd206e32f01e),
    .INIT_65(256'h022ffd206bd0982f022ffd0bc3a2f01e022ffd206e501001022ffd207132b20f),
    .INIT_66(256'h022ffd2070d01102022ffd2071b010a0022ffd250000b203022ffd206e319801),
    .INIT_67(256'h022ffd0bc0603f03022ffd206ef208eb022ffd206ef208be022ffd206e5208db),
    .INIT_68(256'h022ffd0bc042ff0f022ffd206bd2fe0e022ffd0bc052fd0d022ffd206bd2fc0c),
    .INIT_69(256'h022ffd207290bf0f022ffd207f00be0e022ffd206e30bd0d022ffd206bd0bc0c),
    .INIT_6A(256'h022ffd0d504208f5022ffd09502208db022ffd206e501100022ffd2070501020),
    .INIT_6B(256'h022ffd09c1c22017022ffd227c6361b1022ffd208020d001022ffd3a7af0b001),
    .INIT_6C(256'h022ffd0bb0220918022ffd09f1f208ca022ffd09e1e208b2022ffd09d1d221b4),
    .INIT_6D(256'h022ffd13d001f000022ffd10cb00b017022ffd14b061d000022ffd14b060b016),
    .INIT_6E(256'h022ffd2fe361f000022ffd2ff3b0b019022ffd13f001f000022ffd13e000b018),
    .INIT_6F(256'h022ffd206bd1f000022ffd0bc3b0b01b022ffd2fc341f000022ffd2fd350b01a),
    .INIT_70(256'h022ffd206bd1f000022ffd0bc350b01d022ffd206bd1f000022ffd0bc360b01c),
    .INIT_71(256'h022ffd20707324d4022ffd206e31d002022ffd206bd0b032022ffd0bc34361d0),
    .INIT_72(256'h022ffd3a7ce208ac022ffd0d5042f03a022ffd206e511001022ffd207050b03a),
    .INIT_73(256'h022ffd0bd3522008022ffd0bc3432481022ffd227e41d001022ffd208020b032),
    .INIT_74(256'h022ffd01b001d800022ffd01a0430901022ffd0bf3b0d001022ffd0be360b001),
    .INIT_75(256'h022ffd2062f0b017022ffd09f072f034022ffd2062f0b016022ffd2068132206),
    .INIT_76(256'h022ffd2062f0b019022ffd09d072f036022ffd2062f0b018022ffd09e072f035),
    .INIT_77(256'h022ffd206bd0b01b022ffd00cd02f03c022ffd206bd0b01a022ffd09c072f03b),
    .INIT_78(256'h022ffd206bd0b01d022ffd00cf02f03e022ffd206bd0b01c022ffd00ce02f03d),
    .INIT_79(256'h022ffd206e5208ca022ffd20719208b2022ffd20707208f8022ffd206e32f03f),
    .INIT_7A(256'h022ffd14c001c010022ffd0d5040b134022ffd01c000b016022ffd206ef20918),
    .INIT_7B(256'h022ffd250000b018022ffd206e31e010022ffd206bd0b135022ffd11c010b017),
    .INIT_7C(256'h022ffd2b80c0b13b022ffd206e50b019022ffd207271e010022ffd207290b136),
    .INIT_7D(256'h022ffd2b02c1e010022ffd206bd0b13c022ffd09c0c0b01a022ffd2b03c1e010),
    .INIT_7E(256'h022ffd09c0c0b01c022ffd2b01c1e010022ffd206bd0b13d022ffd09c0c0b01b),
    .INIT_7F(256'h022ffd206bd0b13f022ffd09c0c0b01d022ffd2b00c1e010022ffd206bd0b13e),
    .INITP_00(256'hea15a290fa6fe877d9dba57d72cca12d14b159ababa08b319c592e80886e0692),
    .INITP_01(256'ha4b8a8fea4bd9ae7cddb60df043aace77efafe20a3b95bfa6e5bb0943dfa4470),
    .INITP_02(256'hf25f61e05b6fe2d3e16174d0e14b7fe3e9e9f27ed451d33306331b0c1c851020),
    .INITP_03(256'h415b696ad0ec63664d5e5153f57f47c9eedf7febf96873c0e6c5c3fef8c9cdd7),
    .INITP_04(256'h65f8eee0f7c5c15ef4e2556d70f953f46267e8d473fef3d977ebe766624be7e7),
    .INITP_05(256'h4f6175c965cd7afe5e4cdcfad0e04e6ce0ce69794e6840655f6743d65ae147e0),
    .INITP_06(256'h5e69e4eddbd55f50c65c59517f6968f95becf86ac06fca7355f9cecb7951eb6d),
    .INITP_07(256'h5ffa5c7246fbdce7def2447259f1d87c487243f6527352727cf15f7852eac253),
    .INITP_08(256'he7f8f57060ea61f6676f7b61f4eafe77e66f796175ea7ff6ecfe7f656065dde1),
    .INITP_09(256'hffdaea7dfedde96acbea78f67464e7f665f879f77a7c79eafff6686460f07ff8),
    .INITP_0A(256'h73e95667f74ecd714cee4c65f0705d756ed0dde04277536c6df1c869facb7cef),
    .INITP_0B(256'h5573647b57c06fd172edd843eed4efff7a7159e9c963fee8d6ed6bc643747343),
    .INITP_0C(256'he262e567d641e76ad7627fc2456ce1f359716fdece4c49f7766745e8df7c65e3),
    .INITP_0D(256'hda7e71c14e79efc04bcf7863434d7bf1c57cd8d4e0c0f149c1556cc7ee4f7fc4),
    .INITP_0E(256'hd052535ff27e71fff65f75534b7e754ad870795ae67169445f69de67da67da65),
    .INITP_0F(256'hd1c95c524ac254ca43d749ddecf7d85661e45351467b63ed6d424ffad3c85050),
