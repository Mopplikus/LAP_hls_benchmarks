	component kernel_2mm is
		port (
			clock                : in  std_logic                     := 'X';             -- clk
			resetn               : in  std_logic                     := 'X';             -- reset_n
			start                : in  std_logic                     := 'X';             -- valid
			busy                 : out std_logic;                                        -- stall
			done                 : out std_logic;                                        -- valid
			stall                : in  std_logic                     := 'X';             -- stall
			alpha                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			beta                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			A                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			B                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			C                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			D                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			avmm_0_rw_address    : out std_logic_vector(63 downto 0);                    -- address
			avmm_0_rw_byteenable : out std_logic_vector(7 downto 0);                     -- byteenable
			avmm_0_rw_read       : out std_logic;                                        -- read
			avmm_0_rw_readdata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			avmm_0_rw_write      : out std_logic;                                        -- write
			avmm_0_rw_writedata  : out std_logic_vector(63 downto 0)                     -- writedata
		);
	end component kernel_2mm;

	u0 : component kernel_2mm
		port map (
			clock                => CONNECTED_TO_clock,                --     clock.clk
			resetn               => CONNECTED_TO_resetn,               --     reset.reset_n
			start                => CONNECTED_TO_start,                --      call.valid
			busy                 => CONNECTED_TO_busy,                 --          .stall
			done                 => CONNECTED_TO_done,                 --    return.valid
			stall                => CONNECTED_TO_stall,                --          .stall
			alpha                => CONNECTED_TO_alpha,                --     alpha.data
			beta                 => CONNECTED_TO_beta,                 --      beta.data
			A                    => CONNECTED_TO_A,                    --         A.data
			B                    => CONNECTED_TO_B,                    --         B.data
			C                    => CONNECTED_TO_C,                    --         C.data
			D                    => CONNECTED_TO_D,                    --         D.data
			avmm_0_rw_address    => CONNECTED_TO_avmm_0_rw_address,    -- avmm_0_rw.address
			avmm_0_rw_byteenable => CONNECTED_TO_avmm_0_rw_byteenable, --          .byteenable
			avmm_0_rw_read       => CONNECTED_TO_avmm_0_rw_read,       --          .read
			avmm_0_rw_readdata   => CONNECTED_TO_avmm_0_rw_readdata,   --          .readdata
			avmm_0_rw_write      => CONNECTED_TO_avmm_0_rw_write,      --          .write
			avmm_0_rw_writedata  => CONNECTED_TO_avmm_0_rw_writedata   --          .writedata
		);

